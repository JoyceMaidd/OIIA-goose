reg [2:0] frame3 [0:24][0:24] = '{
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd1,3'd5,3'd5,3'd1,3'd1,3'd1,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd1,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd2,3'd2,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd1,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd2,3'd1,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd1,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd4,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd5,3'd5,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
    '{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}
};