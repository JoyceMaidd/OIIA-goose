// frame0.svh — 25x25 goose sprite ROM
reg [2:0] frame0 [0:24][0:24];

initial begin
    frame0[0][0] = 4'd0;
    frame0[0][1] = 4'd0;
    frame0[0][2] = 4'd0;
    frame0[0][3] = 4'd0;
    frame0[0][4] = 4'd0;
    frame0[0][5] = 4'd0;
    frame0[0][6] = 4'd0;
    frame0[0][7] = 4'd0;
    frame0[0][8] = 4'd0;
    frame0[0][9] = 4'd0;
    frame0[0][10] = 4'd0;
    frame0[0][11] = 4'd0;
    frame0[0][12] = 4'd0;
    frame0[0][13] = 4'd0;
    frame0[0][14] = 4'd0;
    frame0[0][15] = 4'd0;
    frame0[0][16] = 4'd0;
    frame0[0][17] = 4'd0;
    frame0[0][18] = 4'd0;
    frame0[0][19] = 4'd0;
    frame0[0][20] = 4'd0;
    frame0[0][21] = 4'd0;
    frame0[0][22] = 4'd0;
    frame0[0][23] = 4'd0;
    frame0[0][24] = 4'd0;
    frame0[1][0] = 4'd0;
    frame0[1][1] = 4'd0;
    frame0[1][2] = 4'd0;
    frame0[1][3] = 4'd0;
    frame0[1][4] = 4'd0;
    frame0[1][5] = 4'd0;
    frame0[1][6] = 4'd0;
    frame0[1][7] = 4'd0;
    frame0[1][8] = 4'd0;
    frame0[1][9] = 4'd0;
    frame0[1][10] = 4'd1;
    frame0[1][11] = 4'd1;
    frame0[1][12] = 4'd1;
    frame0[1][13] = 4'd1;
    frame0[1][14] = 4'd1;
    frame0[1][15] = 4'd0;
    frame0[1][16] = 4'd0;
    frame0[1][17] = 4'd0;
    frame0[1][18] = 4'd0;
    frame0[1][19] = 4'd0;
    frame0[1][20] = 4'd0;
    frame0[1][21] = 4'd0;
    frame0[1][22] = 4'd0;
    frame0[1][23] = 4'd0;
    frame0[1][24] = 4'd0;
    frame0[2][0] = 4'd0;
    frame0[2][1] = 4'd0;
    frame0[2][2] = 4'd0;
    frame0[2][3] = 4'd0;
    frame0[2][4] = 4'd0;
    frame0[2][5] = 4'd0;
    frame0[2][6] = 4'd0;
    frame0[2][7] = 4'd0;
    frame0[2][8] = 4'd0;
    frame0[2][9] = 4'd2;
    frame0[2][10] = 4'd2;
    frame0[2][11] = 4'd2;
    frame0[2][12] = 4'd2;
    frame0[2][13] = 4'd2;
    frame0[2][14] = 4'd2;
    frame0[2][15] = 4'd2;
    frame0[2][16] = 4'd0;
    frame0[2][17] = 4'd0;
    frame0[2][18] = 4'd0;
    frame0[2][19] = 4'd0;
    frame0[2][20] = 4'd0;
    frame0[2][21] = 4'd0;
    frame0[2][22] = 4'd0;
    frame0[2][23] = 4'd0;
    frame0[2][24] = 4'd0;
    frame0[3][0] = 4'd0;
    frame0[3][1] = 4'd0;
    frame0[3][2] = 4'd0;
    frame0[3][3] = 4'd0;
    frame0[3][4] = 4'd0;
    frame0[3][5] = 4'd0;
    frame0[3][6] = 4'd0;
    frame0[3][7] = 4'd0;
    frame0[3][8] = 4'd0;
    frame0[3][9] = 4'd1;
    frame0[3][10] = 4'd1;
    frame0[3][11] = 4'd2;
    frame0[3][12] = 4'd2;
    frame0[3][13] = 4'd2;
    frame0[3][14] = 4'd1;
    frame0[3][15] = 4'd1;
    frame0[3][16] = 4'd0;
    frame0[3][17] = 4'd0;
    frame0[3][18] = 4'd0;
    frame0[3][19] = 4'd0;
    frame0[3][20] = 4'd0;
    frame0[3][21] = 4'd0;
    frame0[3][22] = 4'd0;
    frame0[3][23] = 4'd0;
    frame0[3][24] = 4'd0;
    frame0[4][0] = 4'd0;
    frame0[4][1] = 4'd0;
    frame0[4][2] = 4'd0;
    frame0[4][3] = 4'd0;
    frame0[4][4] = 4'd0;
    frame0[4][5] = 4'd0;
    frame0[4][6] = 4'd0;
    frame0[4][7] = 4'd0;
    frame0[4][8] = 4'd0;
    frame0[4][9] = 4'd3;
    frame0[4][10] = 4'd1;
    frame0[4][11] = 4'd2;
    frame0[4][12] = 4'd2;
    frame0[4][13] = 4'd2;
    frame0[4][14] = 4'd1;
    frame0[4][15] = 4'd3;
    frame0[4][16] = 4'd0;
    frame0[4][17] = 4'd0;
    frame0[4][18] = 4'd0;
    frame0[4][19] = 4'd0;
    frame0[4][20] = 4'd0;
    frame0[4][21] = 4'd0;
    frame0[4][22] = 4'd0;
    frame0[4][23] = 4'd0;
    frame0[4][24] = 4'd0;
    frame0[5][0] = 4'd0;
    frame0[5][1] = 4'd0;
    frame0[5][2] = 4'd0;
    frame0[5][3] = 4'd0;
    frame0[5][4] = 4'd0;
    frame0[5][5] = 4'd0;
    frame0[5][6] = 4'd0;
    frame0[5][7] = 4'd0;
    frame0[5][8] = 4'd0;
    frame0[5][9] = 4'd1;
    frame0[5][10] = 4'd1;
    frame0[5][11] = 4'd3;
    frame0[5][12] = 4'd1;
    frame0[5][13] = 4'd3;
    frame0[5][14] = 4'd1;
    frame0[5][15] = 4'd1;
    frame0[5][16] = 4'd0;
    frame0[5][17] = 4'd0;
    frame0[5][18] = 4'd0;
    frame0[5][19] = 4'd0;
    frame0[5][20] = 4'd0;
    frame0[5][21] = 4'd0;
    frame0[5][22] = 4'd0;
    frame0[5][23] = 4'd0;
    frame0[5][24] = 4'd0;
    frame0[6][0] = 4'd0;
    frame0[6][1] = 4'd0;
    frame0[6][2] = 4'd0;
    frame0[6][3] = 4'd0;
    frame0[6][4] = 4'd0;
    frame0[6][5] = 4'd0;
    frame0[6][6] = 4'd0;
    frame0[6][7] = 4'd0;
    frame0[6][8] = 4'd0;
    frame0[6][9] = 4'd0;
    frame0[6][10] = 4'd0;
    frame0[6][11] = 4'd1;
    frame0[6][12] = 4'd1;
    frame0[6][13] = 4'd1;
    frame0[6][14] = 4'd0;
    frame0[6][15] = 4'd0;
    frame0[6][16] = 4'd0;
    frame0[6][17] = 4'd0;
    frame0[6][18] = 4'd0;
    frame0[6][19] = 4'd0;
    frame0[6][20] = 4'd0;
    frame0[6][21] = 4'd0;
    frame0[6][22] = 4'd0;
    frame0[6][23] = 4'd0;
    frame0[6][24] = 4'd0;
    frame0[7][0] = 4'd0;
    frame0[7][1] = 4'd0;
    frame0[7][2] = 4'd0;
    frame0[7][3] = 4'd0;
    frame0[7][4] = 4'd0;
    frame0[7][5] = 4'd0;
    frame0[7][6] = 4'd0;
    frame0[7][7] = 4'd0;
    frame0[7][8] = 4'd0;
    frame0[7][9] = 4'd0;
    frame0[7][10] = 4'd0;
    frame0[7][11] = 4'd1;
    frame0[7][12] = 4'd2;
    frame0[7][13] = 4'd1;
    frame0[7][14] = 4'd0;
    frame0[7][15] = 4'd0;
    frame0[7][16] = 4'd0;
    frame0[7][17] = 4'd0;
    frame0[7][18] = 4'd0;
    frame0[7][19] = 4'd0;
    frame0[7][20] = 4'd0;
    frame0[7][21] = 4'd0;
    frame0[7][22] = 4'd0;
    frame0[7][23] = 4'd0;
    frame0[7][24] = 4'd0;
    frame0[8][0] = 4'd0;
    frame0[8][1] = 4'd0;
    frame0[8][2] = 4'd0;
    frame0[8][3] = 4'd0;
    frame0[8][4] = 4'd0;
    frame0[8][5] = 4'd0;
    frame0[8][6] = 4'd0;
    frame0[8][7] = 4'd0;
    frame0[8][8] = 4'd0;
    frame0[8][9] = 4'd0;
    frame0[8][10] = 4'd0;
    frame0[8][11] = 4'd1;
    frame0[8][12] = 4'd2;
    frame0[8][13] = 4'd1;
    frame0[8][14] = 4'd0;
    frame0[8][15] = 4'd0;
    frame0[8][16] = 4'd0;
    frame0[8][17] = 4'd0;
    frame0[8][18] = 4'd0;
    frame0[8][19] = 4'd0;
    frame0[8][20] = 4'd0;
    frame0[8][21] = 4'd0;
    frame0[8][22] = 4'd0;
    frame0[8][23] = 4'd0;
    frame0[8][24] = 4'd0;
    frame0[9][0] = 4'd0;
    frame0[9][1] = 4'd0;
    frame0[9][2] = 4'd0;
    frame0[9][3] = 4'd0;
    frame0[9][4] = 4'd0;
    frame0[9][5] = 4'd0;
    frame0[9][6] = 4'd0;
    frame0[9][7] = 4'd0;
    frame0[9][8] = 4'd0;
    frame0[9][9] = 4'd0;
    frame0[9][10] = 4'd0;
    frame0[9][11] = 4'd1;
    frame0[9][12] = 4'd2;
    frame0[9][13] = 4'd1;
    frame0[9][14] = 4'd0;
    frame0[9][15] = 4'd0;
    frame0[9][16] = 4'd0;
    frame0[9][17] = 4'd0;
    frame0[9][18] = 4'd0;
    frame0[9][19] = 4'd0;
    frame0[9][20] = 4'd0;
    frame0[9][21] = 4'd0;
    frame0[9][22] = 4'd0;
    frame0[9][23] = 4'd0;
    frame0[9][24] = 4'd0;
    frame0[10][0] = 4'd0;
    frame0[10][1] = 4'd0;
    frame0[10][2] = 4'd0;
    frame0[10][3] = 4'd0;
    frame0[10][4] = 4'd0;
    frame0[10][5] = 4'd0;
    frame0[10][6] = 4'd0;
    frame0[10][7] = 4'd0;
    frame0[10][8] = 4'd0;
    frame0[10][9] = 4'd0;
    frame0[10][10] = 4'd1;
    frame0[10][11] = 4'd1;
    frame0[10][12] = 4'd2;
    frame0[10][13] = 4'd1;
    frame0[10][14] = 4'd1;
    frame0[10][15] = 4'd0;
    frame0[10][16] = 4'd0;
    frame0[10][17] = 4'd0;
    frame0[10][18] = 4'd0;
    frame0[10][19] = 4'd0;
    frame0[10][20] = 4'd0;
    frame0[10][21] = 4'd0;
    frame0[10][22] = 4'd0;
    frame0[10][23] = 4'd0;
    frame0[10][24] = 4'd0;
    frame0[11][0] = 4'd0;
    frame0[11][1] = 4'd0;
    frame0[11][2] = 4'd0;
    frame0[11][3] = 4'd0;
    frame0[11][4] = 4'd0;
    frame0[11][5] = 4'd0;
    frame0[11][6] = 4'd0;
    frame0[11][7] = 4'd0;
    frame0[11][8] = 4'd0;
    frame0[11][9] = 4'd1;
    frame0[11][10] = 4'd2;
    frame0[11][11] = 4'd4;
    frame0[11][12] = 4'd4;
    frame0[11][13] = 4'd4;
    frame0[11][14] = 4'd2;
    frame0[11][15] = 4'd1;
    frame0[11][16] = 4'd0;
    frame0[11][17] = 4'd0;
    frame0[11][18] = 4'd0;
    frame0[11][19] = 4'd0;
    frame0[11][20] = 4'd0;
    frame0[11][21] = 4'd0;
    frame0[11][22] = 4'd0;
    frame0[11][23] = 4'd0;
    frame0[11][24] = 4'd0;
    frame0[12][0] = 4'd0;
    frame0[12][1] = 4'd0;
    frame0[12][2] = 4'd0;
    frame0[12][3] = 4'd0;
    frame0[12][4] = 4'd0;
    frame0[12][5] = 4'd0;
    frame0[12][6] = 4'd0;
    frame0[12][7] = 4'd0;
    frame0[12][8] = 4'd0;
    frame0[12][9] = 4'd2;
    frame0[12][10] = 4'd2;
    frame0[12][11] = 4'd4;
    frame0[12][12] = 4'd4;
    frame0[12][13] = 4'd4;
    frame0[12][14] = 4'd2;
    frame0[12][15] = 4'd2;
    frame0[12][16] = 4'd0;
    frame0[12][17] = 4'd0;
    frame0[12][18] = 4'd0;
    frame0[12][19] = 4'd0;
    frame0[12][20] = 4'd0;
    frame0[12][21] = 4'd0;
    frame0[12][22] = 4'd0;
    frame0[12][23] = 4'd0;
    frame0[12][24] = 4'd0;
    frame0[13][0] = 4'd0;
    frame0[13][1] = 4'd0;
    frame0[13][2] = 4'd0;
    frame0[13][3] = 4'd0;
    frame0[13][4] = 4'd0;
    frame0[13][5] = 4'd0;
    frame0[13][6] = 4'd1;
    frame0[13][7] = 4'd1;
    frame0[13][8] = 4'd2;
    frame0[13][9] = 4'd4;
    frame0[13][10] = 4'd4;
    frame0[13][11] = 4'd4;
    frame0[13][12] = 4'd4;
    frame0[13][13] = 4'd4;
    frame0[13][14] = 4'd4;
    frame0[13][15] = 4'd4;
    frame0[13][16] = 4'd2;
    frame0[13][17] = 4'd1;
    frame0[13][18] = 4'd1;
    frame0[13][19] = 4'd0;
    frame0[13][20] = 4'd0;
    frame0[13][21] = 4'd0;
    frame0[13][22] = 4'd0;
    frame0[13][23] = 4'd0;
    frame0[13][24] = 4'd0;
    frame0[14][0] = 4'd0;
    frame0[14][1] = 4'd0;
    frame0[14][2] = 4'd0;
    frame0[14][3] = 4'd0;
    frame0[14][4] = 4'd0;
    frame0[14][5] = 4'd1;
    frame0[14][6] = 4'd1;
    frame0[14][7] = 4'd2;
    frame0[14][8] = 4'd2;
    frame0[14][9] = 4'd4;
    frame0[14][10] = 4'd4;
    frame0[14][11] = 4'd4;
    frame0[14][12] = 4'd4;
    frame0[14][13] = 4'd4;
    frame0[14][14] = 4'd4;
    frame0[14][15] = 4'd4;
    frame0[14][16] = 4'd2;
    frame0[14][17] = 4'd2;
    frame0[14][18] = 4'd1;
    frame0[14][19] = 4'd1;
    frame0[14][20] = 4'd0;
    frame0[14][21] = 4'd0;
    frame0[14][22] = 4'd0;
    frame0[14][23] = 4'd0;
    frame0[14][24] = 4'd0;
    frame0[15][0] = 4'd0;
    frame0[15][1] = 4'd0;
    frame0[15][2] = 4'd0;
    frame0[15][3] = 4'd0;
    frame0[15][4] = 4'd0;
    frame0[15][5] = 4'd1;
    frame0[15][6] = 4'd2;
    frame0[15][7] = 4'd2;
    frame0[15][8] = 4'd2;
    frame0[15][9] = 4'd4;
    frame0[15][10] = 4'd4;
    frame0[15][11] = 4'd4;
    frame0[15][12] = 4'd4;
    frame0[15][13] = 4'd4;
    frame0[15][14] = 4'd4;
    frame0[15][15] = 4'd4;
    frame0[15][16] = 4'd2;
    frame0[15][17] = 4'd2;
    frame0[15][18] = 4'd2;
    frame0[15][19] = 4'd1;
    frame0[15][20] = 4'd0;
    frame0[15][21] = 4'd0;
    frame0[15][22] = 4'd0;
    frame0[15][23] = 4'd0;
    frame0[15][24] = 4'd0;
    frame0[16][0] = 4'd0;
    frame0[16][1] = 4'd0;
    frame0[16][2] = 4'd0;
    frame0[16][3] = 4'd0;
    frame0[16][4] = 4'd0;
    frame0[16][5] = 4'd1;
    frame0[16][6] = 4'd1;
    frame0[16][7] = 4'd2;
    frame0[16][8] = 4'd1;
    frame0[16][9] = 4'd5;
    frame0[16][10] = 4'd4;
    frame0[16][11] = 4'd4;
    frame0[16][12] = 4'd4;
    frame0[16][13] = 4'd4;
    frame0[16][14] = 4'd4;
    frame0[16][15] = 4'd5;
    frame0[16][16] = 4'd1;
    frame0[16][17] = 4'd2;
    frame0[16][18] = 4'd1;
    frame0[16][19] = 4'd1;
    frame0[16][20] = 4'd0;
    frame0[16][21] = 4'd0;
    frame0[16][22] = 4'd0;
    frame0[16][23] = 4'd0;
    frame0[16][24] = 4'd0;
    frame0[17][0] = 4'd0;
    frame0[17][1] = 4'd0;
    frame0[17][2] = 4'd0;
    frame0[17][3] = 4'd0;
    frame0[17][4] = 4'd0;
    frame0[17][5] = 4'd0;
    frame0[17][6] = 4'd1;
    frame0[17][7] = 4'd1;
    frame0[17][8] = 4'd1;
    frame0[17][9] = 4'd2;
    frame0[17][10] = 4'd5;
    frame0[17][11] = 4'd4;
    frame0[17][12] = 4'd4;
    frame0[17][13] = 4'd4;
    frame0[17][14] = 4'd5;
    frame0[17][15] = 4'd2;
    frame0[17][16] = 4'd1;
    frame0[17][17] = 4'd1;
    frame0[17][18] = 4'd1;
    frame0[17][19] = 4'd0;
    frame0[17][20] = 4'd0;
    frame0[17][21] = 4'd0;
    frame0[17][22] = 4'd0;
    frame0[17][23] = 4'd0;
    frame0[17][24] = 4'd0;
    frame0[18][0] = 4'd0;
    frame0[18][1] = 4'd0;
    frame0[18][2] = 4'd0;
    frame0[18][3] = 4'd0;
    frame0[18][4] = 4'd0;
    frame0[18][5] = 4'd0;
    frame0[18][6] = 4'd0;
    frame0[18][7] = 4'd1;
    frame0[18][8] = 4'd1;
    frame0[18][9] = 4'd2;
    frame0[18][10] = 4'd2;
    frame0[18][11] = 4'd5;
    frame0[18][12] = 4'd5;
    frame0[18][13] = 4'd5;
    frame0[18][14] = 4'd2;
    frame0[18][15] = 4'd2;
    frame0[18][16] = 4'd1;
    frame0[18][17] = 4'd1;
    frame0[18][18] = 4'd0;
    frame0[18][19] = 4'd0;
    frame0[18][20] = 4'd0;
    frame0[18][21] = 4'd0;
    frame0[18][22] = 4'd0;
    frame0[18][23] = 4'd0;
    frame0[18][24] = 4'd0;
    frame0[19][0] = 4'd0;
    frame0[19][1] = 4'd0;
    frame0[19][2] = 4'd0;
    frame0[19][3] = 4'd0;
    frame0[19][4] = 4'd0;
    frame0[19][5] = 4'd0;
    frame0[19][6] = 4'd0;
    frame0[19][7] = 4'd0;
    frame0[19][8] = 4'd0;
    frame0[19][9] = 4'd1;
    frame0[19][10] = 4'd2;
    frame0[19][11] = 4'd2;
    frame0[19][12] = 4'd5;
    frame0[19][13] = 4'd2;
    frame0[19][14] = 4'd2;
    frame0[19][15] = 4'd1;
    frame0[19][16] = 4'd0;
    frame0[19][17] = 4'd0;
    frame0[19][18] = 4'd0;
    frame0[19][19] = 4'd0;
    frame0[19][20] = 4'd0;
    frame0[19][21] = 4'd0;
    frame0[19][22] = 4'd0;
    frame0[19][23] = 4'd0;
    frame0[19][24] = 4'd0;
    frame0[20][0] = 4'd0;
    frame0[20][1] = 4'd0;
    frame0[20][2] = 4'd0;
    frame0[20][3] = 4'd0;
    frame0[20][4] = 4'd0;
    frame0[20][5] = 4'd0;
    frame0[20][6] = 4'd0;
    frame0[20][7] = 4'd0;
    frame0[20][8] = 4'd0;
    frame0[20][9] = 4'd1;
    frame0[20][10] = 4'd0;
    frame0[20][11] = 4'd1;
    frame0[20][12] = 4'd2;
    frame0[20][13] = 4'd1;
    frame0[20][14] = 4'd0;
    frame0[20][15] = 4'd1;
    frame0[20][16] = 4'd0;
    frame0[20][17] = 4'd0;
    frame0[20][18] = 4'd0;
    frame0[20][19] = 4'd0;
    frame0[20][20] = 4'd0;
    frame0[20][21] = 4'd0;
    frame0[20][22] = 4'd0;
    frame0[20][23] = 4'd0;
    frame0[20][24] = 4'd0;
    frame0[21][0] = 4'd0;
    frame0[21][1] = 4'd0;
    frame0[21][2] = 4'd0;
    frame0[21][3] = 4'd0;
    frame0[21][4] = 4'd0;
    frame0[21][5] = 4'd0;
    frame0[21][6] = 4'd0;
    frame0[21][7] = 4'd0;
    frame0[21][8] = 4'd0;
    frame0[21][9] = 4'd1;
    frame0[21][10] = 4'd0;
    frame0[21][11] = 4'd0;
    frame0[21][12] = 4'd1;
    frame0[21][13] = 4'd0;
    frame0[21][14] = 4'd0;
    frame0[21][15] = 4'd1;
    frame0[21][16] = 4'd0;
    frame0[21][17] = 4'd0;
    frame0[21][18] = 4'd0;
    frame0[21][19] = 4'd0;
    frame0[21][20] = 4'd0;
    frame0[21][21] = 4'd0;
    frame0[21][22] = 4'd0;
    frame0[21][23] = 4'd0;
    frame0[21][24] = 4'd0;
    frame0[22][0] = 4'd0;
    frame0[22][1] = 4'd0;
    frame0[22][2] = 4'd0;
    frame0[22][3] = 4'd0;
    frame0[22][4] = 4'd0;
    frame0[22][5] = 4'd0;
    frame0[22][6] = 4'd0;
    frame0[22][7] = 4'd0;
    frame0[22][8] = 4'd0;
    frame0[22][9] = 4'd1;
    frame0[22][10] = 4'd0;
    frame0[22][11] = 4'd0;
    frame0[22][12] = 4'd0;
    frame0[22][13] = 4'd0;
    frame0[22][14] = 4'd0;
    frame0[22][15] = 4'd1;
    frame0[22][16] = 4'd0;
    frame0[22][17] = 4'd0;
    frame0[22][18] = 4'd0;
    frame0[22][19] = 4'd0;
    frame0[22][20] = 4'd0;
    frame0[22][21] = 4'd0;
    frame0[22][22] = 4'd0;
    frame0[22][23] = 4'd0;
    frame0[22][24] = 4'd0;
    frame0[23][0] = 4'd0;
    frame0[23][1] = 4'd0;
    frame0[23][2] = 4'd0;
    frame0[23][3] = 4'd0;
    frame0[23][4] = 4'd0;
    frame0[23][5] = 4'd0;
    frame0[23][6] = 4'd0;
    frame0[23][7] = 4'd0;
    frame0[23][8] = 4'd0;
    frame0[23][9] = 4'd1;
    frame0[23][10] = 4'd1;
    frame0[23][11] = 4'd0;
    frame0[23][12] = 4'd0;
    frame0[23][13] = 4'd0;
    frame0[23][14] = 4'd1;
    frame0[23][15] = 4'd1;
    frame0[23][16] = 4'd0;
    frame0[23][17] = 4'd0;
    frame0[23][18] = 4'd0;
    frame0[23][19] = 4'd0;
    frame0[23][20] = 4'd0;
    frame0[23][21] = 4'd0;
    frame0[23][22] = 4'd0;
    frame0[23][23] = 4'd0;
    frame0[23][24] = 4'd0;
    frame0[24][0] = 4'd0;
    frame0[24][1] = 4'd0;
    frame0[24][2] = 4'd0;
    frame0[24][3] = 4'd0;
    frame0[24][4] = 4'd0;
    frame0[24][5] = 4'd0;
    frame0[24][6] = 4'd0;
    frame0[24][7] = 4'd0;
    frame0[24][8] = 4'd1;
    frame0[24][9] = 4'd1;
    frame0[24][10] = 4'd0;
    frame0[24][11] = 4'd1;
    frame0[24][12] = 4'd0;
    frame0[24][13] = 4'd1;
    frame0[24][14] = 4'd0;
    frame0[24][15] = 4'd1;
    frame0[24][16] = 4'd1;
    frame0[24][17] = 4'd0;
    frame0[24][18] = 4'd0;
    frame0[24][19] = 4'd0;
    frame0[24][20] = 4'd0;
    frame0[24][21] = 4'd0;
    frame0[24][22] = 4'd0;
    frame0[24][23] = 4'd0;
    frame0[24][24] = 4'd0;
end
