reg [5:0] frame2[7:0][31:0];
initial begin
    frame2[0][0] = 6'd0;
    frame2[1][0] = 6'd0;
    frame2[2][0] = 6'd0;
    frame2[3][0] = 6'd0;
    frame2[4][0] = 6'd0;
    frame2[5][0] = 6'd0;
    frame2[6][0] = 6'd0;
    frame2[7][0] = 6'd0;
    frame2[0][1] = 6'd0;
    frame2[1][1] = 6'd0;
    frame2[2][1] = 6'd0;
    frame2[3][1] = 6'd0;
    frame2[4][1] = 6'd0;
    frame2[5][1] = 6'd0;
    frame2[6][1] = 6'd0;
    frame2[7][1] = 6'd0;
    frame2[0][2] = 6'd0;
    frame2[1][2] = 6'd0;
    frame2[2][2] = 6'd0;
    frame2[3][2] = 6'd7;
    frame2[4][2] = 6'd8;
    frame2[5][2] = 6'd0;
    frame2[6][2] = 6'd0;
    frame2[7][2] = 6'd0;
    frame2[0][3] = 6'd0;
    frame2[1][3] = 6'd0;
    frame2[2][3] = 6'd0;
    frame2[3][3] = 6'd5;
    frame2[4][3] = 6'd4;
    frame2[5][3] = 6'd0;
    frame2[6][3] = 6'd0;
    frame2[7][3] = 6'd0;
    frame2[0][4] = 6'd0;
    frame2[1][4] = 6'd0;
    frame2[2][4] = 6'd0;
    frame2[3][4] = 6'd5;
    frame2[4][4] = 6'd4;
    frame2[5][4] = 6'd0;
    frame2[6][4] = 6'd0;
    frame2[7][4] = 6'd0;
    frame2[0][5] = 6'd0;
    frame2[1][5] = 6'd0;
    frame2[2][5] = 6'd0;
    frame2[3][5] = 6'd22;
    frame2[4][5] = 6'd33;
    frame2[5][5] = 6'd0;
    frame2[6][5] = 6'd0;
    frame2[7][5] = 6'd0;
    frame2[0][6] = 6'd0;
    frame2[1][6] = 6'd0;
    frame2[2][6] = 6'd0;
    frame2[3][6] = 6'd39;
    frame2[4][6] = 6'd60;
    frame2[5][6] = 6'd0;
    frame2[6][6] = 6'd0;
    frame2[7][6] = 6'd0;
    frame2[0][7] = 6'd0;
    frame2[1][7] = 6'd0;
    frame2[2][7] = 6'd0;
    frame2[3][7] = 6'd3;
    frame2[4][7] = 6'd2;
    frame2[5][7] = 6'd0;
    frame2[6][7] = 6'd0;
    frame2[7][7] = 6'd0;
    frame2[0][8] = 6'd0;
    frame2[1][8] = 6'd0;
    frame2[2][8] = 6'd0;
    frame2[3][8] = 6'd3;
    frame2[4][8] = 6'd2;
    frame2[5][8] = 6'd0;
    frame2[6][8] = 6'd0;
    frame2[7][8] = 6'd0;
    frame2[0][9] = 6'd0;
    frame2[1][9] = 6'd0;
    frame2[2][9] = 6'd0;
    frame2[3][9] = 6'd3;
    frame2[4][9] = 6'd2;
    frame2[5][9] = 6'd0;
    frame2[6][9] = 6'd0;
    frame2[7][9] = 6'd0;
    frame2[0][10] = 6'd0;
    frame2[1][10] = 6'd0;
    frame2[2][10] = 6'd0;
    frame2[3][10] = 6'd3;
    frame2[4][10] = 6'd2;
    frame2[5][10] = 6'd0;
    frame2[6][10] = 6'd0;
    frame2[7][10] = 6'd0;
    frame2[0][11] = 6'd0;
    frame2[1][11] = 6'd0;
    frame2[2][11] = 6'd0;
    frame2[3][11] = 6'd3;
    frame2[4][11] = 6'd2;
    frame2[5][11] = 6'd0;
    frame2[6][11] = 6'd0;
    frame2[7][11] = 6'd0;
    frame2[0][12] = 6'd0;
    frame2[1][12] = 6'd0;
    frame2[2][12] = 6'd0;
    frame2[3][12] = 6'd3;
    frame2[4][12] = 6'd2;
    frame2[5][12] = 6'd0;
    frame2[6][12] = 6'd0;
    frame2[7][12] = 6'd0;
    frame2[0][13] = 6'd0;
    frame2[1][13] = 6'd0;
    frame2[2][13] = 6'd0;
    frame2[3][13] = 6'd3;
    frame2[4][13] = 6'd2;
    frame2[5][13] = 6'd0;
    frame2[6][13] = 6'd0;
    frame2[7][13] = 6'd0;
    frame2[0][14] = 6'd0;
    frame2[1][14] = 6'd0;
    frame2[2][14] = 6'd0;
    frame2[3][14] = 6'd5;
    frame2[4][14] = 6'd4;
    frame2[5][14] = 6'd0;
    frame2[6][14] = 6'd0;
    frame2[7][14] = 6'd0;
    frame2[0][15] = 6'd0;
    frame2[1][15] = 6'd0;
    frame2[2][15] = 6'd0;
    frame2[3][15] = 6'd1;
    frame2[4][15] = 6'd1;
    frame2[5][15] = 6'd0;
    frame2[6][15] = 6'd0;
    frame2[7][15] = 6'd0;
    frame2[0][16] = 6'd0;
    frame2[1][16] = 6'd0;
    frame2[2][16] = 6'd3;
    frame2[3][16] = 6'd1;
    frame2[4][16] = 6'd1;
    frame2[5][16] = 6'd2;
    frame2[6][16] = 6'd0;
    frame2[7][16] = 6'd0;
    frame2[0][17] = 6'd0;
    frame2[1][17] = 6'd0;
    frame2[2][17] = 6'd7;
    frame2[3][17] = 6'd1;
    frame2[4][17] = 6'd1;
    frame2[5][17] = 6'd8;
    frame2[6][17] = 6'd0;
    frame2[7][17] = 6'd0;
    frame2[0][18] = 6'd0;
    frame2[1][18] = 6'd0;
    frame2[2][18] = 6'd5;
    frame2[3][18] = 6'd1;
    frame2[4][18] = 6'd1;
    frame2[5][18] = 6'd4;
    frame2[6][18] = 6'd0;
    frame2[7][18] = 6'd0;
    frame2[0][19] = 6'd0;
    frame2[1][19] = 6'd0;
    frame2[2][19] = 6'd1;
    frame2[3][19] = 6'd1;
    frame2[4][19] = 6'd1;
    frame2[5][19] = 6'd1;
    frame2[6][19] = 6'd0;
    frame2[7][19] = 6'd0;
    frame2[0][20] = 6'd0;
    frame2[1][20] = 6'd0;
    frame2[2][20] = 6'd5;
    frame2[3][20] = 6'd1;
    frame2[4][20] = 6'd1;
    frame2[5][20] = 6'd4;
    frame2[6][20] = 6'd0;
    frame2[7][20] = 6'd0;
    frame2[0][21] = 6'd0;
    frame2[1][21] = 6'd0;
    frame2[2][21] = 6'd0;
    frame2[3][21] = 6'd1;
    frame2[4][21] = 6'd1;
    frame2[5][21] = 6'd0;
    frame2[6][21] = 6'd0;
    frame2[7][21] = 6'd0;
    frame2[0][22] = 6'd0;
    frame2[1][22] = 6'd0;
    frame2[2][22] = 6'd30;
    frame2[3][22] = 6'd5;
    frame2[4][22] = 6'd4;
    frame2[5][22] = 6'd23;
    frame2[6][22] = 6'd0;
    frame2[7][22] = 6'd0;
    frame2[0][23] = 6'd0;
    frame2[1][23] = 6'd0;
    frame2[2][23] = 6'd28;
    frame2[3][23] = 6'd3;
    frame2[4][23] = 6'd2;
    frame2[5][23] = 6'd24;
    frame2[6][23] = 6'd0;
    frame2[7][23] = 6'd0;
    frame2[0][24] = 6'd0;
    frame2[1][24] = 6'd0;
    frame2[2][24] = 6'd16;
    frame2[3][24] = 6'd56;
    frame2[4][24] = 6'd36;
    frame2[5][24] = 6'd11;
    frame2[6][24] = 6'd0;
    frame2[7][24] = 6'd0;
    frame2[0][25] = 6'd0;
    frame2[1][25] = 6'd0;
    frame2[2][25] = 6'd0;
    frame2[3][25] = 6'd30;
    frame2[4][25] = 6'd23;
    frame2[5][25] = 6'd0;
    frame2[6][25] = 6'd0;
    frame2[7][25] = 6'd0;
    frame2[0][26] = 6'd0;
    frame2[1][26] = 6'd0;
    frame2[2][26] = 6'd0;
    frame2[3][26] = 6'd28;
    frame2[4][26] = 6'd24;
    frame2[5][26] = 6'd0;
    frame2[6][26] = 6'd0;
    frame2[7][26] = 6'd0;
    frame2[0][27] = 6'd0;
    frame2[1][27] = 6'd0;
    frame2[2][27] = 6'd0;
    frame2[3][27] = 6'd0;
    frame2[4][27] = 6'd0;
    frame2[5][27] = 6'd0;
    frame2[6][27] = 6'd0;
    frame2[7][27] = 6'd0;
    frame2[0][28] = 6'd0;
    frame2[1][28] = 6'd0;
    frame2[2][28] = 6'd0;
    frame2[3][28] = 6'd0;
    frame2[4][28] = 6'd0;
    frame2[5][28] = 6'd0;
    frame2[6][28] = 6'd0;
    frame2[7][28] = 6'd0;
    frame2[0][29] = 6'd0;
    frame2[1][29] = 6'd0;
    frame2[2][29] = 6'd0;
    frame2[3][29] = 6'd0;
    frame2[4][29] = 6'd0;
    frame2[5][29] = 6'd0;
    frame2[6][29] = 6'd0;
    frame2[7][29] = 6'd0;
    frame2[0][30] = 6'd0;
    frame2[1][30] = 6'd0;
    frame2[2][30] = 6'd0;
    frame2[3][30] = 6'd0;
    frame2[4][30] = 6'd0;
    frame2[5][30] = 6'd0;
    frame2[6][30] = 6'd0;
    frame2[7][30] = 6'd0;
    frame2[0][31] = 6'd0;
    frame2[1][31] = 6'd0;
    frame2[2][31] = 6'd0;
    frame2[3][31] = 6'd0;
    frame2[4][31] = 6'd0;
    frame2[5][31] = 6'd0;
    frame2[6][31] = 6'd0;
    frame2[7][31] = 6'd0;
end
