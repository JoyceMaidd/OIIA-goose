reg [5:0] frame0[7:0][31:0];
initial begin
    frame0[0][0] = 6'd0;
    frame0[1][0] = 6'd0;
    frame0[2][0] = 6'd0;
    frame0[3][0] = 6'd0;
    frame0[4][0] = 6'd0;
    frame0[5][0] = 6'd0;
    frame0[6][0] = 6'd0;
    frame0[7][0] = 6'd0;
    frame0[0][1] = 6'd0;
    frame0[1][1] = 6'd0;
    frame0[2][1] = 6'd0;
    frame0[3][1] = 6'd0;
    frame0[4][1] = 6'd0;
    frame0[5][1] = 6'd0;
    frame0[6][1] = 6'd0;
    frame0[7][1] = 6'd0;
    frame0[0][2] = 6'd0;
    frame0[1][2] = 6'd0;
    frame0[2][2] = 6'd0;
    frame0[3][2] = 6'd7;
    frame0[4][2] = 6'd8;
    frame0[5][2] = 6'd0;
    frame0[6][2] = 6'd0;
    frame0[7][2] = 6'd0;
    frame0[0][3] = 6'd0;
    frame0[1][3] = 6'd0;
    frame0[2][3] = 6'd0;
    frame0[3][3] = 6'd1;
    frame0[4][3] = 6'd1;
    frame0[5][3] = 6'd0;
    frame0[6][3] = 6'd0;
    frame0[7][3] = 6'd0;
    frame0[0][4] = 6'd0;
    frame0[1][4] = 6'd0;
    frame0[2][4] = 6'd0;
    frame0[3][4] = 6'd7;
    frame0[4][4] = 6'd8;
    frame0[5][4] = 6'd0;
    frame0[6][4] = 6'd0;
    frame0[7][4] = 6'd0;
    frame0[0][5] = 6'd0;
    frame0[1][5] = 6'd0;
    frame0[2][5] = 6'd0;
    frame0[3][5] = 6'd53;
    frame0[4][5] = 6'd44;
    frame0[5][5] = 6'd0;
    frame0[6][5] = 6'd0;
    frame0[7][5] = 6'd0;
    frame0[0][6] = 6'd0;
    frame0[1][6] = 6'd0;
    frame0[2][6] = 6'd0;
    frame0[3][6] = 6'd58;
    frame0[4][6] = 6'd51;
    frame0[5][6] = 6'd0;
    frame0[6][6] = 6'd0;
    frame0[7][6] = 6'd0;
    frame0[0][7] = 6'd0;
    frame0[1][7] = 6'd0;
    frame0[2][7] = 6'd0;
    frame0[3][7] = 6'd32;
    frame0[4][7] = 6'd27;
    frame0[5][7] = 6'd0;
    frame0[6][7] = 6'd0;
    frame0[7][7] = 6'd0;
    frame0[0][8] = 6'd0;
    frame0[1][8] = 6'd0;
    frame0[2][8] = 6'd0;
    frame0[3][8] = 6'd0;
    frame0[4][8] = 6'd0;
    frame0[5][8] = 6'd0;
    frame0[6][8] = 6'd0;
    frame0[7][8] = 6'd0;
    frame0[0][9] = 6'd0;
    frame0[1][9] = 6'd0;
    frame0[2][9] = 6'd0;
    frame0[3][9] = 6'd3;
    frame0[4][9] = 6'd2;
    frame0[5][9] = 6'd0;
    frame0[6][9] = 6'd0;
    frame0[7][9] = 6'd0;
    frame0[0][10] = 6'd0;
    frame0[1][10] = 6'd0;
    frame0[2][10] = 6'd0;
    frame0[3][10] = 6'd3;
    frame0[4][10] = 6'd2;
    frame0[5][10] = 6'd0;
    frame0[6][10] = 6'd0;
    frame0[7][10] = 6'd0;
    frame0[0][11] = 6'd0;
    frame0[1][11] = 6'd0;
    frame0[2][11] = 6'd0;
    frame0[3][11] = 6'd3;
    frame0[4][11] = 6'd2;
    frame0[5][11] = 6'd0;
    frame0[6][11] = 6'd0;
    frame0[7][11] = 6'd0;
    frame0[0][12] = 6'd0;
    frame0[1][12] = 6'd0;
    frame0[2][12] = 6'd0;
    frame0[3][12] = 6'd3;
    frame0[4][12] = 6'd2;
    frame0[5][12] = 6'd0;
    frame0[6][12] = 6'd0;
    frame0[7][12] = 6'd0;
    frame0[0][13] = 6'd0;
    frame0[1][13] = 6'd0;
    frame0[2][13] = 6'd0;
    frame0[3][13] = 6'd3;
    frame0[4][13] = 6'd2;
    frame0[5][13] = 6'd0;
    frame0[6][13] = 6'd0;
    frame0[7][13] = 6'd0;
    frame0[0][14] = 6'd0;
    frame0[1][14] = 6'd0;
    frame0[2][14] = 6'd0;
    frame0[3][14] = 6'd45;
    frame0[4][14] = 6'd46;
    frame0[5][14] = 6'd0;
    frame0[6][14] = 6'd0;
    frame0[7][14] = 6'd0;
    frame0[0][15] = 6'd0;
    frame0[1][15] = 6'd0;
    frame0[2][15] = 6'd0;
    frame0[3][15] = 6'd14;
    frame0[4][15] = 6'd12;
    frame0[5][15] = 6'd0;
    frame0[6][15] = 6'd0;
    frame0[7][15] = 6'd0;
    frame0[0][16] = 6'd0;
    frame0[1][16] = 6'd0;
    frame0[2][16] = 6'd3;
    frame0[3][16] = 6'd17;
    frame0[4][16] = 6'd15;
    frame0[5][16] = 6'd2;
    frame0[6][16] = 6'd0;
    frame0[7][16] = 6'd0;
    frame0[0][17] = 6'd0;
    frame0[1][17] = 6'd0;
    frame0[2][17] = 6'd7;
    frame0[3][17] = 6'd6;
    frame0[4][17] = 6'd6;
    frame0[5][17] = 6'd8;
    frame0[6][17] = 6'd0;
    frame0[7][17] = 6'd0;
    frame0[0][18] = 6'd0;
    frame0[1][18] = 6'd0;
    frame0[2][18] = 6'd5;
    frame0[3][18] = 6'd6;
    frame0[4][18] = 6'd6;
    frame0[5][18] = 6'd4;
    frame0[6][18] = 6'd0;
    frame0[7][18] = 6'd0;
    frame0[0][19] = 6'd0;
    frame0[1][19] = 6'd0;
    frame0[2][19] = 6'd1;
    frame0[3][19] = 6'd6;
    frame0[4][19] = 6'd6;
    frame0[5][19] = 6'd1;
    frame0[6][19] = 6'd0;
    frame0[7][19] = 6'd0;
    frame0[0][20] = 6'd0;
    frame0[1][20] = 6'd0;
    frame0[2][20] = 6'd18;
    frame0[3][20] = 6'd6;
    frame0[4][20] = 6'd6;
    frame0[5][20] = 6'd19;
    frame0[6][20] = 6'd0;
    frame0[7][20] = 6'd0;
    frame0[0][21] = 6'd0;
    frame0[1][21] = 6'd0;
    frame0[2][21] = 6'd43;
    frame0[3][21] = 6'd17;
    frame0[4][21] = 6'd15;
    frame0[5][21] = 6'd48;
    frame0[6][21] = 6'd0;
    frame0[7][21] = 6'd0;
    frame0[0][22] = 6'd0;
    frame0[1][22] = 6'd0;
    frame0[2][22] = 6'd3;
    frame0[3][22] = 6'd14;
    frame0[4][22] = 6'd12;
    frame0[5][22] = 6'd2;
    frame0[6][22] = 6'd0;
    frame0[7][22] = 6'd0;
    frame0[0][23] = 6'd0;
    frame0[1][23] = 6'd0;
    frame0[2][23] = 6'd0;
    frame0[3][23] = 6'd1;
    frame0[4][23] = 6'd1;
    frame0[5][23] = 6'd0;
    frame0[6][23] = 6'd0;
    frame0[7][23] = 6'd0;
    frame0[0][24] = 6'd0;
    frame0[1][24] = 6'd0;
    frame0[2][24] = 6'd0;
    frame0[3][24] = 6'd5;
    frame0[4][24] = 6'd4;
    frame0[5][24] = 6'd0;
    frame0[6][24] = 6'd0;
    frame0[7][24] = 6'd0;
    frame0[0][25] = 6'd0;
    frame0[1][25] = 6'd0;
    frame0[2][25] = 6'd0;
    frame0[3][25] = 6'd7;
    frame0[4][25] = 6'd8;
    frame0[5][25] = 6'd0;
    frame0[6][25] = 6'd0;
    frame0[7][25] = 6'd0;
    frame0[0][26] = 6'd0;
    frame0[1][26] = 6'd0;
    frame0[2][26] = 6'd0;
    frame0[3][26] = 6'd3;
    frame0[4][26] = 6'd2;
    frame0[5][26] = 6'd0;
    frame0[6][26] = 6'd0;
    frame0[7][26] = 6'd0;
    frame0[0][27] = 6'd0;
    frame0[1][27] = 6'd0;
    frame0[2][27] = 6'd0;
    frame0[3][27] = 6'd0;
    frame0[4][27] = 6'd0;
    frame0[5][27] = 6'd0;
    frame0[6][27] = 6'd0;
    frame0[7][27] = 6'd0;
    frame0[0][28] = 6'd0;
    frame0[1][28] = 6'd0;
    frame0[2][28] = 6'd0;
    frame0[3][28] = 6'd0;
    frame0[4][28] = 6'd0;
    frame0[5][28] = 6'd0;
    frame0[6][28] = 6'd0;
    frame0[7][28] = 6'd0;
    frame0[0][29] = 6'd0;
    frame0[1][29] = 6'd0;
    frame0[2][29] = 6'd0;
    frame0[3][29] = 6'd0;
    frame0[4][29] = 6'd0;
    frame0[5][29] = 6'd0;
    frame0[6][29] = 6'd0;
    frame0[7][29] = 6'd0;
    frame0[0][30] = 6'd0;
    frame0[1][30] = 6'd0;
    frame0[2][30] = 6'd0;
    frame0[3][30] = 6'd0;
    frame0[4][30] = 6'd0;
    frame0[5][30] = 6'd0;
    frame0[6][30] = 6'd0;
    frame0[7][30] = 6'd0;
    frame0[0][31] = 6'd0;
    frame0[1][31] = 6'd0;
    frame0[2][31] = 6'd0;
    frame0[3][31] = 6'd0;
    frame0[4][31] = 6'd0;
    frame0[5][31] = 6'd0;
    frame0[6][31] = 6'd0;
    frame0[7][31] = 6'd0;
end
