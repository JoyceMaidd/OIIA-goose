reg [2:0] frame3 [0:1][0:1];

initial begin
    frame3[0][0] = 3'h0;
    frame3[0][1] = 3'h0;
    // frame3[0][2] = 3'h0;
    // frame3[0][3] = 3'h0;
    // frame3[0][4] = 3'h0;
    // frame3[0][5] = 3'h0;
    // frame3[0][6] = 3'h0;
    // frame3[0][7] = 3'h0;
    // frame3[0][8] = 3'h0;
    // frame3[0][9] = 3'h0;
    // frame3[0][10] = 3'h0;
    // frame3[0][11] = 3'h0;
    // frame3[0][12] = 3'h0;
    // frame3[0][13] = 3'h0;
    // frame3[0][14] = 3'h0;
    // frame3[0][15] = 3'h0;
    // frame3[0][16] = 3'h0;
    // frame3[0][17] = 3'h0;
    // frame3[0][18] = 3'h0;
    // frame3[0][19] = 3'h0;
    // frame3[0][20] = 3'h0;
    // frame3[0][21] = 3'h0;
    // frame3[0][22] = 3'h0;
    // frame3[0][23] = 3'h0;
    // frame3[0][24] = 3'h0;
    // frame3[0][25] = 3'h0;
    // frame3[0][26] = 3'h0;
    // frame3[0][27] = 3'h0;
    // frame3[0][28] = 3'h0;
    // frame3[0][29] = 3'h0;
    // frame3[0][30] = 3'h0;
    // frame3[0][31] = 3'h0;
    frame3[1][0] = 3'h0;
    frame3[1][1] = 3'h0;
    // frame3[1][2] = 3'h0;
    // frame3[1][3] = 3'h0;
    // frame3[1][4] = 3'h0;
    // frame3[1][5] = 3'h0;
    // frame3[1][6] = 3'h0;
    // frame3[1][7] = 3'h0;
    // frame3[1][8] = 3'h0;
    // frame3[1][9] = 3'h0;
    // frame3[1][10] = 3'h0;
    // frame3[1][11] = 3'h0;
    // frame3[1][12] = 3'h0;
    // frame3[1][13] = 3'h0;
    // frame3[1][14] = 3'h0;
    // frame3[1][15] = 3'h0;
    // frame3[1][16] = 3'h0;
    // frame3[1][17] = 3'h0;
    // frame3[1][18] = 3'h0;
    // frame3[1][19] = 3'h0;
    // frame3[1][20] = 3'h1;
    // frame3[1][21] = 3'h1;
    // frame3[1][22] = 3'h1;
    // frame3[1][23] = 3'h1;
    // frame3[1][24] = 3'h1;
    // frame3[1][25] = 3'h1;
    // frame3[1][26] = 3'h0;
    // frame3[1][27] = 3'h0;
    // frame3[1][28] = 3'h0;
    // frame3[1][29] = 3'h0;
    // frame3[1][30] = 3'h0;
    // frame3[1][31] = 3'h0;
    // frame3[2][0] = 3'h0;
    // frame3[2][1] = 3'h0;
    // frame3[2][2] = 3'h0;
    // frame3[2][3] = 3'h0;
    // frame3[2][4] = 3'h0;
    // frame3[2][5] = 3'h0;
    // frame3[2][6] = 3'h0;
    // frame3[2][7] = 3'h0;
    // frame3[2][8] = 3'h0;
    // frame3[2][9] = 3'h0;
    // frame3[2][10] = 3'h0;
    // frame3[2][11] = 3'h0;
    // frame3[2][12] = 3'h0;
    // frame3[2][13] = 3'h0;
    // frame3[2][14] = 3'h0;
    // frame3[2][15] = 3'h0;
    // frame3[2][16] = 3'h0;
    // frame3[2][17] = 3'h0;
    // frame3[2][18] = 3'h0;
    // frame3[2][19] = 3'h1;
    // frame3[2][20] = 3'h1;
    // frame3[2][21] = 3'h2;
    // frame3[2][22] = 3'h2;
    // frame3[2][23] = 3'h2;
    // frame3[2][24] = 3'h2;
    // frame3[2][25] = 3'h1;
    // frame3[2][26] = 3'h1;
    // frame3[2][27] = 3'h0;
    // frame3[2][28] = 3'h0;
    // frame3[2][29] = 3'h0;
    // frame3[2][30] = 3'h0;
    // frame3[2][31] = 3'h0;
    // frame3[3][0] = 3'h0;
    // frame3[3][1] = 3'h0;
    // frame3[3][2] = 3'h0;
    // frame3[3][3] = 3'h0;
    // frame3[3][4] = 3'h0;
    // frame3[3][5] = 3'h0;
    // frame3[3][6] = 3'h0;
    // frame3[3][7] = 3'h0;
    // frame3[3][8] = 3'h0;
    // frame3[3][9] = 3'h0;
    // frame3[3][10] = 3'h0;
    // frame3[3][11] = 3'h0;
    // frame3[3][12] = 3'h0;
    // frame3[3][13] = 3'h0;
    // frame3[3][14] = 3'h0;
    // frame3[3][15] = 3'h0;
    // frame3[3][16] = 3'h0;
    // frame3[3][17] = 3'h0;
    // frame3[3][18] = 3'h0;
    // frame3[3][19] = 3'h1;
    // frame3[3][20] = 3'h2;
    // frame3[3][21] = 3'h2;
    // frame3[3][22] = 3'h2;
    // frame3[3][23] = 3'h2;
    // frame3[3][24] = 3'h2;
    // frame3[3][25] = 3'h2;
    // frame3[3][26] = 3'h1;
    // frame3[3][27] = 3'h1;
    // frame3[3][28] = 3'h0;
    // frame3[3][29] = 3'h0;
    // frame3[3][30] = 3'h0;
    // frame3[3][31] = 3'h0;
    // frame3[4][0] = 3'h0;
    // frame3[4][1] = 3'h0;
    // frame3[4][2] = 3'h0;
    // frame3[4][3] = 3'h0;
    // frame3[4][4] = 3'h0;
    // frame3[4][5] = 3'h0;
    // frame3[4][6] = 3'h0;
    // frame3[4][7] = 3'h0;
    // frame3[4][8] = 3'h0;
    // frame3[4][9] = 3'h0;
    // frame3[4][10] = 3'h0;
    // frame3[4][11] = 3'h0;
    // frame3[4][12] = 3'h0;
    // frame3[4][13] = 3'h0;
    // frame3[4][14] = 3'h0;
    // frame3[4][15] = 3'h0;
    // frame3[4][16] = 3'h0;
    // frame3[4][17] = 3'h0;
    // frame3[4][18] = 3'h0;
    // frame3[4][19] = 3'h1;
    // frame3[4][20] = 3'h2;
    // frame3[4][21] = 3'h2;
    // frame3[4][22] = 3'h2;
    // frame3[4][23] = 3'h1;
    // frame3[4][24] = 3'h1;
    // frame3[4][25] = 3'h2;
    // frame3[4][26] = 3'h2;
    // frame3[4][27] = 3'h1;
    // frame3[4][28] = 3'h0;
    // frame3[4][29] = 3'h0;
    // frame3[4][30] = 3'h0;
    // frame3[4][31] = 3'h0;
    // frame3[5][0] = 3'h0;
    // frame3[5][1] = 3'h0;
    // frame3[5][2] = 3'h0;
    // frame3[5][3] = 3'h0;
    // frame3[5][4] = 3'h0;
    // frame3[5][5] = 3'h0;
    // frame3[5][6] = 3'h0;
    // frame3[5][7] = 3'h0;
    // frame3[5][8] = 3'h0;
    // frame3[5][9] = 3'h0;
    // frame3[5][10] = 3'h0;
    // frame3[5][11] = 3'h0;
    // frame3[5][12] = 3'h0;
    // frame3[5][13] = 3'h0;
    // frame3[5][14] = 3'h0;
    // frame3[5][15] = 3'h0;
    // frame3[5][16] = 3'h0;
    // frame3[5][17] = 3'h0;
    // frame3[5][18] = 3'h0;
    // frame3[5][19] = 3'h1;
    // frame3[5][20] = 3'h2;
    // frame3[5][21] = 3'h2;
    // frame3[5][22] = 3'h2;
    // frame3[5][23] = 3'h2;
    // frame3[5][24] = 3'h1;
    // frame3[5][25] = 3'h2;
    // frame3[5][26] = 3'h2;
    // frame3[5][27] = 3'h1;
    // frame3[5][28] = 3'h0;
    // frame3[5][29] = 3'h0;
    // frame3[5][30] = 3'h0;
    // frame3[5][31] = 3'h0;
    // frame3[6][0] = 3'h0;
    // frame3[6][1] = 3'h0;
    // frame3[6][2] = 3'h0;
    // frame3[6][3] = 3'h0;
    // frame3[6][4] = 3'h0;
    // frame3[6][5] = 3'h0;
    // frame3[6][6] = 3'h0;
    // frame3[6][7] = 3'h0;
    // frame3[6][8] = 3'h0;
    // frame3[6][9] = 3'h0;
    // frame3[6][10] = 3'h0;
    // frame3[6][11] = 3'h0;
    // frame3[6][12] = 3'h0;
    // frame3[6][13] = 3'h0;
    // frame3[6][14] = 3'h0;
    // frame3[6][15] = 3'h0;
    // frame3[6][16] = 3'h0;
    // frame3[6][17] = 3'h0;
    // frame3[6][18] = 3'h0;
    // frame3[6][19] = 3'h1;
    // frame3[6][20] = 3'h3;
    // frame3[6][21] = 3'h2;
    // frame3[6][22] = 3'h2;
    // frame3[6][23] = 3'h2;
    // frame3[6][24] = 3'h2;
    // frame3[6][25] = 3'h2;
    // frame3[6][26] = 3'h2;
    // frame3[6][27] = 3'h1;
    // frame3[6][28] = 3'h1;
    // frame3[6][29] = 3'h1;
    // frame3[6][30] = 3'h1;
    // frame3[6][31] = 3'h0;
    // frame3[7][0] = 3'h0;
    // frame3[7][1] = 3'h0;
    // frame3[7][2] = 3'h0;
    // frame3[7][3] = 3'h0;
    // frame3[7][4] = 3'h0;
    // frame3[7][5] = 3'h0;
    // frame3[7][6] = 3'h0;
    // frame3[7][7] = 3'h0;
    // frame3[7][8] = 3'h0;
    // frame3[7][9] = 3'h0;
    // frame3[7][10] = 3'h0;
    // frame3[7][11] = 3'h0;
    // frame3[7][12] = 3'h0;
    // frame3[7][13] = 3'h0;
    // frame3[7][14] = 3'h0;
    // frame3[7][15] = 3'h0;
    // frame3[7][16] = 3'h0;
    // frame3[7][17] = 3'h0;
    // frame3[7][18] = 3'h0;
    // frame3[7][19] = 3'h1;
    // frame3[7][20] = 3'h3;
    // frame3[7][21] = 3'h3;
    // frame3[7][22] = 3'h2;
    // frame3[7][23] = 3'h2;
    // frame3[7][24] = 3'h2;
    // frame3[7][25] = 3'h2;
    // frame3[7][26] = 3'h1;
    // frame3[7][27] = 3'h1;
    // frame3[7][28] = 3'h1;
    // frame3[7][29] = 3'h1;
    // frame3[7][30] = 3'h1;
    // frame3[7][31] = 3'h0;
    // frame3[8][0] = 3'h0;
    // frame3[8][1] = 3'h0;
    // frame3[8][2] = 3'h0;
    // frame3[8][3] = 3'h0;
    // frame3[8][4] = 3'h0;
    // frame3[8][5] = 3'h0;
    // frame3[8][6] = 3'h0;
    // frame3[8][7] = 3'h0;
    // frame3[8][8] = 3'h0;
    // frame3[8][9] = 3'h0;
    // frame3[8][10] = 3'h0;
    // frame3[8][11] = 3'h0;
    // frame3[8][12] = 3'h0;
    // frame3[8][13] = 3'h0;
    // frame3[8][14] = 3'h0;
    // frame3[8][15] = 3'h0;
    // frame3[8][16] = 3'h0;
    // frame3[8][17] = 3'h0;
    // frame3[8][18] = 3'h0;
    // frame3[8][19] = 3'h1;
    // frame3[8][20] = 3'h2;
    // frame3[8][21] = 3'h3;
    // frame3[8][22] = 3'h3;
    // frame3[8][23] = 3'h1;
    // frame3[8][24] = 3'h1;
    // frame3[8][25] = 3'h1;
    // frame3[8][26] = 3'h0;
    // frame3[8][27] = 3'h0;
    // frame3[8][28] = 3'h0;
    // frame3[8][29] = 3'h0;
    // frame3[8][30] = 3'h0;
    // frame3[8][31] = 3'h0;
    // frame3[9][0] = 3'h0;
    // frame3[9][1] = 3'h0;
    // frame3[9][2] = 3'h0;
    // frame3[9][3] = 3'h0;
    // frame3[9][4] = 3'h0;
    // frame3[9][5] = 3'h0;
    // frame3[9][6] = 3'h0;
    // frame3[9][7] = 3'h0;
    // frame3[9][8] = 3'h0;
    // frame3[9][9] = 3'h0;
    // frame3[9][10] = 3'h0;
    // frame3[9][11] = 3'h0;
    // frame3[9][12] = 3'h0;
    // frame3[9][13] = 3'h0;
    // frame3[9][14] = 3'h0;
    // frame3[9][15] = 3'h0;
    // frame3[9][16] = 3'h0;
    // frame3[9][17] = 3'h0;
    // frame3[9][18] = 3'h0;
    // frame3[9][19] = 3'h1;
    // frame3[9][20] = 3'h2;
    // frame3[9][21] = 3'h2;
    // frame3[9][22] = 3'h3;
    // frame3[9][23] = 3'h1;
    // frame3[9][24] = 3'h0;
    // frame3[9][25] = 3'h0;
    // frame3[9][26] = 3'h0;
    // frame3[9][27] = 3'h0;
    // frame3[9][28] = 3'h0;
    // frame3[9][29] = 3'h0;
    // frame3[9][30] = 3'h0;
    // frame3[9][31] = 3'h0;
    // frame3[10][0] = 3'h0;
    // frame3[10][1] = 3'h0;
    // frame3[10][2] = 3'h0;
    // frame3[10][3] = 3'h0;
    // frame3[10][4] = 3'h0;
    // frame3[10][5] = 3'h0;
    // frame3[10][6] = 3'h0;
    // frame3[10][7] = 3'h0;
    // frame3[10][8] = 3'h0;
    // frame3[10][9] = 3'h0;
    // frame3[10][10] = 3'h0;
    // frame3[10][11] = 3'h0;
    // frame3[10][12] = 3'h0;
    // frame3[10][13] = 3'h0;
    // frame3[10][14] = 3'h0;
    // frame3[10][15] = 3'h0;
    // frame3[10][16] = 3'h0;
    // frame3[10][17] = 3'h0;
    // frame3[10][18] = 3'h0;
    // frame3[10][19] = 3'h1;
    // frame3[10][20] = 3'h2;
    // frame3[10][21] = 3'h2;
    // frame3[10][22] = 3'h2;
    // frame3[10][23] = 3'h1;
    // frame3[10][24] = 3'h0;
    // frame3[10][25] = 3'h0;
    // frame3[10][26] = 3'h0;
    // frame3[10][27] = 3'h0;
    // frame3[10][28] = 3'h0;
    // frame3[10][29] = 3'h0;
    // frame3[10][30] = 3'h0;
    // frame3[10][31] = 3'h0;
    // frame3[11][0] = 3'h0;
    // frame3[11][1] = 3'h0;
    // frame3[11][2] = 3'h0;
    // frame3[11][3] = 3'h0;
    // frame3[11][4] = 3'h0;
    // frame3[11][5] = 3'h0;
    // frame3[11][6] = 3'h0;
    // frame3[11][7] = 3'h0;
    // frame3[11][8] = 3'h0;
    // frame3[11][9] = 3'h0;
    // frame3[11][10] = 3'h0;
    // frame3[11][11] = 3'h0;
    // frame3[11][12] = 3'h0;
    // frame3[11][13] = 3'h0;
    // frame3[11][14] = 3'h0;
    // frame3[11][15] = 3'h0;
    // frame3[11][16] = 3'h0;
    // frame3[11][17] = 3'h0;
    // frame3[11][18] = 3'h0;
    // frame3[11][19] = 3'h1;
    // frame3[11][20] = 3'h2;
    // frame3[11][21] = 3'h2;
    // frame3[11][22] = 3'h2;
    // frame3[11][23] = 3'h1;
    // frame3[11][24] = 3'h0;
    // frame3[11][25] = 3'h0;
    // frame3[11][26] = 3'h0;
    // frame3[11][27] = 3'h0;
    // frame3[11][28] = 3'h0;
    // frame3[11][29] = 3'h0;
    // frame3[11][30] = 3'h0;
    // frame3[11][31] = 3'h0;
    // frame3[12][0] = 3'h0;
    // frame3[12][1] = 3'h0;
    // frame3[12][2] = 3'h0;
    // frame3[12][3] = 3'h0;
    // frame3[12][4] = 3'h0;
    // frame3[12][5] = 3'h0;
    // frame3[12][6] = 3'h0;
    // frame3[12][7] = 3'h0;
    // frame3[12][8] = 3'h0;
    // frame3[12][9] = 3'h0;
    // frame3[12][10] = 3'h0;
    // frame3[12][11] = 3'h0;
    // frame3[12][12] = 3'h0;
    // frame3[12][13] = 3'h0;
    // frame3[12][14] = 3'h0;
    // frame3[12][15] = 3'h0;
    // frame3[12][16] = 3'h0;
    // frame3[12][17] = 3'h0;
    // frame3[12][18] = 3'h0;
    // frame3[12][19] = 3'h1;
    // frame3[12][20] = 3'h2;
    // frame3[12][21] = 3'h2;
    // frame3[12][22] = 3'h2;
    // frame3[12][23] = 3'h1;
    // frame3[12][24] = 3'h0;
    // frame3[12][25] = 3'h0;
    // frame3[12][26] = 3'h0;
    // frame3[12][27] = 3'h0;
    // frame3[12][28] = 3'h0;
    // frame3[12][29] = 3'h0;
    // frame3[12][30] = 3'h0;
    // frame3[12][31] = 3'h0;
    // frame3[13][0] = 3'h0;
    // frame3[13][1] = 3'h0;
    // frame3[13][2] = 3'h0;
    // frame3[13][3] = 3'h0;
    // frame3[13][4] = 3'h0;
    // frame3[13][5] = 3'h0;
    // frame3[13][6] = 3'h0;
    // frame3[13][7] = 3'h0;
    // frame3[13][8] = 3'h0;
    // frame3[13][9] = 3'h0;
    // frame3[13][10] = 3'h0;
    // frame3[13][11] = 3'h0;
    // frame3[13][12] = 3'h0;
    // frame3[13][13] = 3'h0;
    // frame3[13][14] = 3'h0;
    // frame3[13][15] = 3'h0;
    // frame3[13][16] = 3'h0;
    // frame3[13][17] = 3'h0;
    // frame3[13][18] = 3'h0;
    // frame3[13][19] = 3'h1;
    // frame3[13][20] = 3'h2;
    // frame3[13][21] = 3'h2;
    // frame3[13][22] = 3'h2;
    // frame3[13][23] = 3'h1;
    // frame3[13][24] = 3'h0;
    // frame3[13][25] = 3'h0;
    // frame3[13][26] = 3'h0;
    // frame3[13][27] = 3'h0;
    // frame3[13][28] = 3'h0;
    // frame3[13][29] = 3'h0;
    // frame3[13][30] = 3'h0;
    // frame3[13][31] = 3'h0;
    // frame3[14][0] = 3'h0;
    // frame3[14][1] = 3'h0;
    // frame3[14][2] = 3'h0;
    // frame3[14][3] = 3'h0;
    // frame3[14][4] = 3'h0;
    // frame3[14][5] = 3'h0;
    // frame3[14][6] = 3'h0;
    // frame3[14][7] = 3'h0;
    // frame3[14][8] = 3'h0;
    // frame3[14][9] = 3'h0;
    // frame3[14][10] = 3'h0;
    // frame3[14][11] = 3'h0;
    // frame3[14][12] = 3'h0;
    // frame3[14][13] = 3'h0;
    // frame3[14][14] = 3'h0;
    // frame3[14][15] = 3'h0;
    // frame3[14][16] = 3'h0;
    // frame3[14][17] = 3'h0;
    // frame3[14][18] = 3'h1;
    // frame3[14][19] = 3'h1;
    // frame3[14][20] = 3'h2;
    // frame3[14][21] = 3'h2;
    // frame3[14][22] = 3'h2;
    // frame3[14][23] = 3'h1;
    // frame3[14][24] = 3'h1;
    // frame3[14][25] = 3'h0;
    // frame3[14][26] = 3'h0;
    // frame3[14][27] = 3'h0;
    // frame3[14][28] = 3'h0;
    // frame3[14][29] = 3'h0;
    // frame3[14][30] = 3'h0;
    // frame3[14][31] = 3'h0;
    // frame3[15][0] = 3'h0;
    // frame3[15][1] = 3'h1;
    // frame3[15][2] = 3'h1;
    // frame3[15][3] = 3'h1;
    // frame3[15][4] = 3'h0;
    // frame3[15][5] = 3'h0;
    // frame3[15][6] = 3'h0;
    // frame3[15][7] = 3'h0;
    // frame3[15][8] = 3'h0;
    // frame3[15][9] = 3'h0;
    // frame3[15][10] = 3'h0;
    // frame3[15][11] = 3'h0;
    // frame3[15][12] = 3'h1;
    // frame3[15][13] = 3'h1;
    // frame3[15][14] = 3'h1;
    // frame3[15][15] = 3'h1;
    // frame3[15][16] = 3'h1;
    // frame3[15][17] = 3'h1;
    // frame3[15][18] = 3'h1;
    // frame3[15][19] = 3'h2;
    // frame3[15][20] = 3'h2;
    // frame3[15][21] = 3'h4;
    // frame3[15][22] = 3'h4;
    // frame3[15][23] = 3'h4;
    // frame3[15][24] = 3'h1;
    // frame3[15][25] = 3'h1;
    // frame3[15][26] = 3'h0;
    // frame3[15][27] = 3'h0;
    // frame3[15][28] = 3'h0;
    // frame3[15][29] = 3'h0;
    // frame3[15][30] = 3'h0;
    // frame3[15][31] = 3'h0;
    // frame3[16][0] = 3'h0;
    // frame3[16][1] = 3'h1;
    // frame3[16][2] = 3'h5;
    // frame3[16][3] = 3'h1;
    // frame3[16][4] = 3'h1;
    // frame3[16][5] = 3'h1;
    // frame3[16][6] = 3'h0;
    // frame3[16][7] = 3'h0;
    // frame3[16][8] = 3'h1;
    // frame3[16][9] = 3'h1;
    // frame3[16][10] = 3'h1;
    // frame3[16][11] = 3'h1;
    // frame3[16][12] = 3'h1;
    // frame3[16][13] = 3'h5;
    // frame3[16][14] = 3'h5;
    // frame3[16][15] = 3'h5;
    // frame3[16][16] = 3'h5;
    // frame3[16][17] = 3'h5;
    // frame3[16][18] = 3'h5;
    // frame3[16][19] = 3'h5;
    // frame3[16][20] = 3'h5;
    // frame3[16][21] = 3'h5;
    // frame3[16][22] = 3'h4;
    // frame3[16][23] = 3'h4;
    // frame3[16][24] = 3'h4;
    // frame3[16][25] = 3'h1;
    // frame3[16][26] = 3'h1;
    // frame3[16][27] = 3'h0;
    // frame3[16][28] = 3'h0;
    // frame3[16][29] = 3'h0;
    // frame3[16][30] = 3'h0;
    // frame3[16][31] = 3'h0;
    // frame3[17][0] = 3'h0;
    // frame3[17][1] = 3'h1;
    // frame3[17][2] = 3'h5;
    // frame3[17][3] = 3'h5;
    // frame3[17][4] = 3'h5;
    // frame3[17][5] = 3'h1;
    // frame3[17][6] = 3'h1;
    // frame3[17][7] = 3'h1;
    // frame3[17][8] = 3'h1;
    // frame3[17][9] = 3'h5;
    // frame3[17][10] = 3'h5;
    // frame3[17][11] = 3'h5;
    // frame3[17][12] = 3'h5;
    // frame3[17][13] = 3'h5;
    // frame3[17][14] = 3'h5;
    // frame3[17][15] = 3'h5;
    // frame3[17][16] = 3'h5;
    // frame3[17][17] = 3'h5;
    // frame3[17][18] = 3'h5;
    // frame3[17][19] = 3'h5;
    // frame3[17][20] = 3'h5;
    // frame3[17][21] = 3'h5;
    // frame3[17][22] = 3'h5;
    // frame3[17][23] = 3'h4;
    // frame3[17][24] = 3'h4;
    // frame3[17][25] = 3'h4;
    // frame3[17][26] = 3'h1;
    // frame3[17][27] = 3'h1;
    // frame3[17][28] = 3'h0;
    // frame3[17][29] = 3'h0;
    // frame3[17][30] = 3'h0;
    // frame3[17][31] = 3'h0;
    // frame3[18][0] = 3'h0;
    // frame3[18][1] = 3'h1;
    // frame3[18][2] = 3'h5;
    // frame3[18][3] = 3'h5;
    // frame3[18][4] = 3'h5;
    // frame3[18][5] = 3'h5;
    // frame3[18][6] = 3'h5;
    // frame3[18][7] = 3'h5;
    // frame3[18][8] = 3'h5;
    // frame3[18][9] = 3'h5;
    // frame3[18][10] = 3'h5;
    // frame3[18][11] = 3'h5;
    // frame3[18][12] = 3'h5;
    // frame3[18][13] = 3'h5;
    // frame3[18][14] = 3'h5;
    // frame3[18][15] = 3'h5;
    // frame3[18][16] = 3'h5;
    // frame3[18][17] = 3'h2;
    // frame3[18][18] = 3'h2;
    // frame3[18][19] = 3'h5;
    // frame3[18][20] = 3'h5;
    // frame3[18][21] = 3'h5;
    // frame3[18][22] = 3'h5;
    // frame3[18][23] = 3'h5;
    // frame3[18][24] = 3'h4;
    // frame3[18][25] = 3'h4;
    // frame3[18][26] = 3'h4;
    // frame3[18][27] = 3'h1;
    // frame3[18][28] = 3'h0;
    // frame3[18][29] = 3'h0;
    // frame3[18][30] = 3'h0;
    // frame3[18][31] = 3'h0;
    // frame3[19][0] = 3'h0;
    // frame3[19][1] = 3'h1;
    // frame3[19][2] = 3'h1;
    // frame3[19][3] = 3'h5;
    // frame3[19][4] = 3'h5;
    // frame3[19][5] = 3'h5;
    // frame3[19][6] = 3'h5;
    // frame3[19][7] = 3'h5;
    // frame3[19][8] = 3'h5;
    // frame3[19][9] = 3'h5;
    // frame3[19][10] = 3'h5;
    // frame3[19][11] = 3'h5;
    // frame3[19][12] = 3'h5;
    // frame3[19][13] = 3'h5;
    // frame3[19][14] = 3'h5;
    // frame3[19][15] = 3'h5;
    // frame3[19][16] = 3'h2;
    // frame3[19][17] = 3'h2;
    // frame3[19][18] = 3'h1;
    // frame3[19][19] = 3'h5;
    // frame3[19][20] = 3'h5;
    // frame3[19][21] = 3'h5;
    // frame3[19][22] = 3'h5;
    // frame3[19][23] = 3'h5;
    // frame3[19][24] = 3'h4;
    // frame3[19][25] = 3'h4;
    // frame3[19][26] = 3'h4;
    // frame3[19][27] = 3'h1;
    // frame3[19][28] = 3'h0;
    // frame3[19][29] = 3'h0;
    // frame3[19][30] = 3'h0;
    // frame3[19][31] = 3'h0;
    // frame3[20][0] = 3'h0;
    // frame3[20][1] = 3'h0;
    // frame3[20][2] = 3'h1;
    // frame3[20][3] = 3'h1;
    // frame3[20][4] = 3'h5;
    // frame3[20][5] = 3'h1;
    // frame3[20][6] = 3'h2;
    // frame3[20][7] = 3'h5;
    // frame3[20][8] = 3'h5;
    // frame3[20][9] = 3'h5;
    // frame3[20][10] = 3'h5;
    // frame3[20][11] = 3'h5;
    // frame3[20][12] = 3'h5;
    // frame3[20][13] = 3'h5;
    // frame3[20][14] = 3'h5;
    // frame3[20][15] = 3'h5;
    // frame3[20][16] = 3'h2;
    // frame3[20][17] = 3'h1;
    // frame3[20][18] = 3'h1;
    // frame3[20][19] = 3'h5;
    // frame3[20][20] = 3'h5;
    // frame3[20][21] = 3'h5;
    // frame3[20][22] = 3'h5;
    // frame3[20][23] = 3'h5;
    // frame3[20][24] = 3'h4;
    // frame3[20][25] = 3'h4;
    // frame3[20][26] = 3'h4;
    // frame3[20][27] = 3'h1;
    // frame3[20][28] = 3'h0;
    // frame3[20][29] = 3'h0;
    // frame3[20][30] = 3'h0;
    // frame3[20][31] = 3'h0;
    // frame3[21][0] = 3'h0;
    // frame3[21][1] = 3'h0;
    // frame3[21][2] = 3'h0;
    // frame3[21][3] = 3'h1;
    // frame3[21][4] = 3'h1;
    // frame3[21][5] = 3'h3;
    // frame3[21][6] = 3'h1;
    // frame3[21][7] = 3'h2;
    // frame3[21][8] = 3'h2;
    // frame3[21][9] = 3'h2;
    // frame3[21][10] = 3'h2;
    // frame3[21][11] = 3'h2;
    // frame3[21][12] = 3'h2;
    // frame3[21][13] = 3'h2;
    // frame3[21][14] = 3'h2;
    // frame3[21][15] = 3'h1;
    // frame3[21][16] = 3'h5;
    // frame3[21][17] = 3'h5;
    // frame3[21][18] = 3'h5;
    // frame3[21][19] = 3'h5;
    // frame3[21][20] = 3'h5;
    // frame3[21][21] = 3'h5;
    // frame3[21][22] = 3'h5;
    // frame3[21][23] = 3'h4;
    // frame3[21][24] = 3'h4;
    // frame3[21][25] = 3'h4;
    // frame3[21][26] = 3'h4;
    // frame3[21][27] = 3'h1;
    // frame3[21][28] = 3'h0;
    // frame3[21][29] = 3'h0;
    // frame3[21][30] = 3'h0;
    // frame3[21][31] = 3'h0;
    // frame3[22][0] = 3'h0;
    // frame3[22][1] = 3'h0;
    // frame3[22][2] = 3'h0;
    // frame3[22][3] = 3'h0;
    // frame3[22][4] = 3'h1;
    // frame3[22][5] = 3'h1;
    // frame3[22][6] = 3'h3;
    // frame3[22][7] = 3'h1;
    // frame3[22][8] = 3'h1;
    // frame3[22][9] = 3'h1;
    // frame3[22][10] = 3'h1;
    // frame3[22][11] = 3'h1;
    // frame3[22][12] = 3'h1;
    // frame3[22][13] = 3'h1;
    // frame3[22][14] = 3'h1;
    // frame3[22][15] = 3'h5;
    // frame3[22][16] = 3'h5;
    // frame3[22][17] = 3'h5;
    // frame3[22][18] = 3'h5;
    // frame3[22][19] = 3'h5;
    // frame3[22][20] = 3'h5;
    // frame3[22][21] = 3'h5;
    // frame3[22][22] = 3'h4;
    // frame3[22][23] = 3'h4;
    // frame3[22][24] = 3'h4;
    // frame3[22][25] = 3'h1;
    // frame3[22][26] = 3'h1;
    // frame3[22][27] = 3'h1;
    // frame3[22][28] = 3'h0;
    // frame3[22][29] = 3'h0;
    // frame3[22][30] = 3'h0;
    // frame3[22][31] = 3'h0;
    // frame3[23][0] = 3'h0;
    // frame3[23][1] = 3'h0;
    // frame3[23][2] = 3'h0;
    // frame3[23][3] = 3'h0;
    // frame3[23][4] = 3'h0;
    // frame3[23][5] = 3'h1;
    // frame3[23][6] = 3'h1;
    // frame3[23][7] = 3'h3;
    // frame3[23][8] = 3'h3;
    // frame3[23][9] = 3'h3;
    // frame3[23][10] = 3'h3;
    // frame3[23][11] = 3'h3;
    // frame3[23][12] = 3'h3;
    // frame3[23][13] = 3'h3;
    // frame3[23][14] = 3'h3;
    // frame3[23][15] = 3'h5;
    // frame3[23][16] = 3'h5;
    // frame3[23][17] = 3'h5;
    // frame3[23][18] = 3'h5;
    // frame3[23][19] = 3'h5;
    // frame3[23][20] = 3'h5;
    // frame3[23][21] = 3'h4;
    // frame3[23][22] = 3'h4;
    // frame3[23][23] = 3'h4;
    // frame3[23][24] = 3'h1;
    // frame3[23][25] = 3'h1;
    // frame3[23][26] = 3'h0;
    // frame3[23][27] = 3'h0;
    // frame3[23][28] = 3'h0;
    // frame3[23][29] = 3'h0;
    // frame3[23][30] = 3'h0;
    // frame3[23][31] = 3'h0;
    // frame3[24][0] = 3'h0;
    // frame3[24][1] = 3'h0;
    // frame3[24][2] = 3'h0;
    // frame3[24][3] = 3'h0;
    // frame3[24][4] = 3'h0;
    // frame3[24][5] = 3'h0;
    // frame3[24][6] = 3'h1;
    // frame3[24][7] = 3'h1;
    // frame3[24][8] = 3'h4;
    // frame3[24][9] = 3'h4;
    // frame3[24][10] = 3'h3;
    // frame3[24][11] = 3'h3;
    // frame3[24][12] = 3'h3;
    // frame3[24][13] = 3'h3;
    // frame3[24][14] = 3'h4;
    // frame3[24][15] = 3'h4;
    // frame3[24][16] = 3'h4;
    // frame3[24][17] = 3'h4;
    // frame3[24][18] = 3'h4;
    // frame3[24][19] = 3'h4;
    // frame3[24][20] = 3'h4;
    // frame3[24][21] = 3'h4;
    // frame3[24][22] = 3'h4;
    // frame3[24][23] = 3'h1;
    // frame3[24][24] = 3'h1;
    // frame3[24][25] = 3'h0;
    // frame3[24][26] = 3'h0;
    // frame3[24][27] = 3'h0;
    // frame3[24][28] = 3'h0;
    // frame3[24][29] = 3'h0;
    // frame3[24][30] = 3'h0;
    // frame3[24][31] = 3'h0;
    // frame3[25][0] = 3'h0;
    // frame3[25][1] = 3'h0;
    // frame3[25][2] = 3'h0;
    // frame3[25][3] = 3'h0;
    // frame3[25][4] = 3'h0;
    // frame3[25][5] = 3'h0;
    // frame3[25][6] = 3'h0;
    // frame3[25][7] = 3'h1;
    // frame3[25][8] = 3'h1;
    // frame3[25][9] = 3'h1;
    // frame3[25][10] = 3'h4;
    // frame3[25][11] = 3'h4;
    // frame3[25][12] = 3'h4;
    // frame3[25][13] = 3'h4;
    // frame3[25][14] = 3'h4;
    // frame3[25][15] = 3'h4;
    // frame3[25][16] = 3'h4;
    // frame3[25][17] = 3'h4;
    // frame3[25][18] = 3'h4;
    // frame3[25][19] = 3'h4;
    // frame3[25][20] = 3'h4;
    // frame3[25][21] = 3'h4;
    // frame3[25][22] = 3'h4;
    // frame3[25][23] = 3'h1;
    // frame3[25][24] = 3'h1;
    // frame3[25][25] = 3'h0;
    // frame3[25][26] = 3'h0;
    // frame3[25][27] = 3'h0;
    // frame3[25][28] = 3'h0;
    // frame3[25][29] = 3'h0;
    // frame3[25][30] = 3'h0;
    // frame3[25][31] = 3'h0;
    // frame3[26][0] = 3'h0;
    // frame3[26][1] = 3'h0;
    // frame3[26][2] = 3'h0;
    // frame3[26][3] = 3'h0;
    // frame3[26][4] = 3'h0;
    // frame3[26][5] = 3'h0;
    // frame3[26][6] = 3'h0;
    // frame3[26][7] = 3'h1;
    // frame3[26][8] = 3'h1;
    // frame3[26][9] = 3'h1;
    // frame3[26][10] = 3'h4;
    // frame3[26][11] = 3'h4;
    // frame3[26][12] = 3'h4;
    // frame3[26][13] = 3'h4;
    // frame3[26][14] = 3'h4;
    // frame3[26][15] = 3'h4;
    // frame3[26][16] = 3'h4;
    // frame3[26][17] = 3'h4;
    // frame3[26][18] = 3'h4;
    // frame3[26][19] = 3'h4;
    // frame3[26][20] = 3'h4;
    // frame3[26][21] = 3'h1;
    // frame3[26][22] = 3'h1;
    // frame3[26][23] = 3'h1;
    // frame3[26][24] = 3'h0;
    // frame3[26][25] = 3'h0;
    // frame3[26][26] = 3'h0;
    // frame3[26][27] = 3'h0;
    // frame3[26][28] = 3'h0;
    // frame3[26][29] = 3'h0;
    // frame3[26][30] = 3'h0;
    // frame3[26][31] = 3'h0;
    // frame3[27][0] = 3'h0;
    // frame3[27][1] = 3'h0;
    // frame3[27][2] = 3'h0;
    // frame3[27][3] = 3'h0;
    // frame3[27][4] = 3'h0;
    // frame3[27][5] = 3'h0;
    // frame3[27][6] = 3'h0;
    // frame3[27][7] = 3'h0;
    // frame3[27][8] = 3'h0;
    // frame3[27][9] = 3'h1;
    // frame3[27][10] = 3'h1;
    // frame3[27][11] = 3'h1;
    // frame3[27][12] = 3'h1;
    // frame3[27][13] = 3'h1;
    // frame3[27][14] = 3'h1;
    // frame3[27][15] = 3'h5;
    // frame3[27][16] = 3'h5;
    // frame3[27][17] = 3'h5;
    // frame3[27][18] = 3'h1;
    // frame3[27][19] = 3'h1;
    // frame3[27][20] = 3'h1;
    // frame3[27][21] = 3'h1;
    // frame3[27][22] = 3'h0;
    // frame3[27][23] = 3'h0;
    // frame3[27][24] = 3'h0;
    // frame3[27][25] = 3'h0;
    // frame3[27][26] = 3'h0;
    // frame3[27][27] = 3'h0;
    // frame3[27][28] = 3'h0;
    // frame3[27][29] = 3'h0;
    // frame3[27][30] = 3'h0;
    // frame3[27][31] = 3'h0;
    // frame3[28][0] = 3'h0;
    // frame3[28][1] = 3'h0;
    // frame3[28][2] = 3'h0;
    // frame3[28][3] = 3'h0;
    // frame3[28][4] = 3'h0;
    // frame3[28][5] = 3'h0;
    // frame3[28][6] = 3'h0;
    // frame3[28][7] = 3'h0;
    // frame3[28][8] = 3'h0;
    // frame3[28][9] = 3'h0;
    // frame3[28][10] = 3'h0;
    // frame3[28][11] = 3'h0;
    // frame3[28][12] = 3'h1;
    // frame3[28][13] = 3'h0;
    // frame3[28][14] = 3'h1;
    // frame3[28][15] = 3'h1;
    // frame3[28][16] = 3'h1;
    // frame3[28][17] = 3'h1;
    // frame3[28][18] = 3'h1;
    // frame3[28][19] = 3'h0;
    // frame3[28][20] = 3'h0;
    // frame3[28][21] = 3'h0;
    // frame3[28][22] = 3'h0;
    // frame3[28][23] = 3'h0;
    // frame3[28][24] = 3'h0;
    // frame3[28][25] = 3'h0;
    // frame3[28][26] = 3'h0;
    // frame3[28][27] = 3'h0;
    // frame3[28][28] = 3'h0;
    // frame3[28][29] = 3'h0;
    // frame3[28][30] = 3'h0;
    // frame3[28][31] = 3'h0;
    // frame3[29][0] = 3'h0;
    // frame3[29][1] = 3'h0;
    // frame3[29][2] = 3'h0;
    // frame3[29][3] = 3'h0;
    // frame3[29][4] = 3'h0;
    // frame3[29][5] = 3'h0;
    // frame3[29][6] = 3'h0;
    // frame3[29][7] = 3'h0;
    // frame3[29][8] = 3'h0;
    // frame3[29][9] = 3'h0;
    // frame3[29][10] = 3'h0;
    // frame3[29][11] = 3'h0;
    // frame3[29][12] = 3'h1;
    // frame3[29][13] = 3'h0;
    // frame3[29][14] = 3'h0;
    // frame3[29][15] = 3'h0;
    // frame3[29][16] = 3'h1;
    // frame3[29][17] = 3'h0;
    // frame3[29][18] = 3'h0;
    // frame3[29][19] = 3'h0;
    // frame3[29][20] = 3'h0;
    // frame3[29][21] = 3'h0;
    // frame3[29][22] = 3'h0;
    // frame3[29][23] = 3'h0;
    // frame3[29][24] = 3'h0;
    // frame3[29][25] = 3'h0;
    // frame3[29][26] = 3'h0;
    // frame3[29][27] = 3'h0;
    // frame3[29][28] = 3'h0;
    // frame3[29][29] = 3'h0;
    // frame3[29][30] = 3'h0;
    // frame3[29][31] = 3'h0;
    // frame3[30][0] = 3'h0;
    // frame3[30][1] = 3'h0;
    // frame3[30][2] = 3'h0;
    // frame3[30][3] = 3'h0;
    // frame3[30][4] = 3'h0;
    // frame3[30][5] = 3'h0;
    // frame3[30][6] = 3'h0;
    // frame3[30][7] = 3'h0;
    // frame3[30][8] = 3'h0;
    // frame3[30][9] = 3'h0;
    // frame3[30][10] = 3'h0;
    // frame3[30][11] = 3'h0;
    // frame3[30][12] = 3'h1;
    // frame3[30][13] = 3'h0;
    // frame3[30][14] = 3'h0;
    // frame3[30][15] = 3'h0;
    // frame3[30][16] = 3'h1;
    // frame3[30][17] = 3'h0;
    // frame3[30][18] = 3'h0;
    // frame3[30][19] = 3'h0;
    // frame3[30][20] = 3'h0;
    // frame3[30][21] = 3'h0;
    // frame3[30][22] = 3'h0;
    // frame3[30][23] = 3'h0;
    // frame3[30][24] = 3'h0;
    // frame3[30][25] = 3'h0;
    // frame3[30][26] = 3'h0;
    // frame3[30][27] = 3'h0;
    // frame3[30][28] = 3'h0;
    // frame3[30][29] = 3'h0;
    // frame3[30][30] = 3'h0;
    // frame3[30][31] = 3'h0;
    // frame3[31][0] = 3'h0;
    // frame3[31][1] = 3'h0;
    // frame3[31][2] = 3'h0;
    // frame3[31][3] = 3'h0;
    // frame3[31][4] = 3'h0;
    // frame3[31][5] = 3'h0;
    // frame3[31][6] = 3'h0;
    // frame3[31][7] = 3'h0;
    // frame3[31][8] = 3'h0;
    // frame3[31][9] = 3'h0;
    // frame3[31][10] = 3'h0;
    // frame3[31][11] = 3'h0;
    // frame3[31][12] = 3'h1;
    // frame3[31][13] = 3'h1;
    // frame3[31][14] = 3'h1;
    // frame3[31][15] = 3'h0;
    // frame3[31][16] = 3'h1;
    // frame3[31][17] = 3'h1;
    // frame3[31][18] = 3'h1;
    // frame3[31][19] = 3'h1;
    // frame3[31][20] = 3'h0;
    // frame3[31][21] = 3'h0;
    // frame3[31][22] = 3'h0;
    // frame3[31][23] = 3'h0;
    // frame3[31][24] = 3'h0;
    // frame3[31][25] = 3'h0;
    // frame3[31][26] = 3'h0;
    // frame3[31][27] = 3'h0;
    // frame3[31][28] = 3'h0;
    // frame3[31][29] = 3'h0;
    // frame3[31][30] = 3'h0;
    // frame3[31][31] = 3'h0;
end
