reg [2:0] frame3 [0:24][0:24];
    initial begin
        frame3[0][0] = 3'd0;
        frame3[0][1] = 3'd0;
        frame3[0][2] = 3'd0;
        frame3[0][3] = 3'd0;
        frame3[0][4] = 3'd0;
        frame3[0][5] = 3'd0;
        frame3[0][6] = 3'd0;
        frame3[0][7] = 3'd0;
        frame3[0][8] = 3'd0;
        frame3[0][9] = 3'd0;
        frame3[0][10] = 3'd0;
        frame3[0][11] = 3'd0;
        frame3[0][12] = 3'd0;
        frame3[0][13] = 3'd0;
        frame3[0][14] = 3'd0;
        frame3[0][15] = 3'd0;
        frame3[0][16] = 3'd0;
        frame3[0][17] = 3'd0;
        frame3[0][18] = 3'd0;
        frame3[0][19] = 3'd0;
        frame3[0][20] = 3'd0;
        frame3[0][21] = 3'd0;
        frame3[0][22] = 3'd0;
        frame3[0][23] = 3'd0;
        frame3[0][24] = 3'd0;
        
        frame3[1][0] = 3'd0;
        frame3[1][1] = 3'd0;
        frame3[1][2] = 3'd0;
        frame3[1][3] = 3'd0;
        frame3[1][4] = 3'd0;
        frame3[1][5] = 3'd0;
        frame3[1][6] = 3'd0;
        frame3[1][7] = 3'd0;
        frame3[1][8] = 3'd0;
        frame3[1][9] = 3'd0;
        frame3[1][10] = 3'd0;
        frame3[1][11] = 3'd0;
        frame3[1][12] = 3'd0;
        frame3[1][13] = 3'd0;
        frame3[1][14] = 3'd0;
        frame3[1][15] = 3'd0;
        frame3[1][16] = 3'd1;
        frame3[1][17] = 3'd1;
        frame3[1][18] = 3'd1;
        frame3[1][19] = 3'd1;
        frame3[1][20] = 3'd0;
        frame3[1][21] = 3'd0;
        frame3[1][22] = 3'd0;
        frame3[1][23] = 3'd0;
        frame3[1][24] = 3'd0;
        
        frame3[2][0] = 3'd0;
        frame3[2][1] = 3'd0;
        frame3[2][2] = 3'd0;
        frame3[2][3] = 3'd0;
        frame3[2][4] = 3'd0;
        frame3[2][5] = 3'd0;
        frame3[2][6] = 3'd0;
        frame3[2][7] = 3'd0;
        frame3[2][8] = 3'd0;
        frame3[2][9] = 3'd0;
        frame3[2][10] = 3'd0;
        frame3[2][11] = 3'd0;
        frame3[2][12] = 3'd0;
        frame3[2][13] = 3'd0;
        frame3[2][14] = 3'd0;
        frame3[2][15] = 3'd1;
        frame3[2][16] = 3'd2;
        frame3[2][17] = 3'd2;
        frame3[2][18] = 3'd2;
        frame3[2][19] = 3'd2;
        frame3[2][20] = 3'd1;
        frame3[2][21] = 3'd1;
        frame3[2][22] = 3'd0;
        frame3[2][23] = 3'd0;
        frame3[2][24] = 3'd0;
        
        frame3[3][0] = 3'd0;
        frame3[3][1] = 3'd0;
        frame3[3][2] = 3'd0;
        frame3[3][3] = 3'd0;
        frame3[3][4] = 3'd0;
        frame3[3][5] = 3'd0;
        frame3[3][6] = 3'd0;
        frame3[3][7] = 3'd0;
        frame3[3][8] = 3'd0;
        frame3[3][9] = 3'd0;
        frame3[3][10] = 3'd0;
        frame3[3][11] = 3'd0;
        frame3[3][12] = 3'd0;
        frame3[3][13] = 3'd0;
        frame3[3][14] = 3'd0;
        frame3[3][15] = 3'd1;
        frame3[3][16] = 3'd2;
        frame3[3][17] = 3'd2;
        frame3[3][18] = 3'd1;
        frame3[3][19] = 3'd1;
        frame3[3][20] = 3'd2;
        frame3[3][21] = 3'd1;
        frame3[3][22] = 3'd0;
        frame3[3][23] = 3'd0;
        frame3[3][24] = 3'd0;
        
        frame3[4][0] = 3'd0;
        frame3[4][1] = 3'd0;
        frame3[4][2] = 3'd0;
        frame3[4][3] = 3'd0;
        frame3[4][4] = 3'd0;
        frame3[4][5] = 3'd0;
        frame3[4][6] = 3'd0;
        frame3[4][7] = 3'd0;
        frame3[4][8] = 3'd0;
        frame3[4][9] = 3'd0;
        frame3[4][10] = 3'd0;
        frame3[4][11] = 3'd0;
        frame3[4][12] = 3'd0;
        frame3[4][13] = 3'd0;
        frame3[4][14] = 3'd0;
        frame3[4][15] = 3'd1;
        frame3[4][16] = 3'd2;
        frame3[4][17] = 3'd2;
        frame3[4][18] = 3'd2;
        frame3[4][19] = 3'd1;
        frame3[4][20] = 3'd2;
        frame3[4][21] = 3'd1;
        frame3[4][22] = 3'd0;
        frame3[4][23] = 3'd0;
        frame3[4][24] = 3'd0;
        
        frame3[5][0] = 3'd0;
        frame3[5][1] = 3'd0;
        frame3[5][2] = 3'd0;
        frame3[5][3] = 3'd0;
        frame3[5][4] = 3'd0;
        frame3[5][5] = 3'd0;
        frame3[5][6] = 3'd0;
        frame3[5][7] = 3'd0;
        frame3[5][8] = 3'd0;
        frame3[5][9] = 3'd0;
        frame3[5][10] = 3'd0;
        frame3[5][11] = 3'd0;
        frame3[5][12] = 3'd0;
        frame3[5][13] = 3'd0;
        frame3[5][14] = 3'd0;
        frame3[5][15] = 3'd1;
        frame3[5][16] = 3'd3;
        frame3[5][17] = 3'd2;
        frame3[5][18] = 3'd2;
        frame3[5][19] = 3'd2;
        frame3[5][20] = 3'd1;
        frame3[5][21] = 3'd1;
        frame3[5][22] = 3'd1;
        frame3[5][23] = 3'd1;
        frame3[5][24] = 3'd0;
        
        frame3[6][0] = 3'd0;
        frame3[6][1] = 3'd0;
        frame3[6][2] = 3'd0;
        frame3[6][3] = 3'd0;
        frame3[6][4] = 3'd0;
        frame3[6][5] = 3'd0;
        frame3[6][6] = 3'd0;
        frame3[6][7] = 3'd0;
        frame3[6][8] = 3'd0;
        frame3[6][9] = 3'd0;
        frame3[6][10] = 3'd0;
        frame3[6][11] = 3'd0;
        frame3[6][12] = 3'd0;
        frame3[6][13] = 3'd0;
        frame3[6][14] = 3'd0;
        frame3[6][15] = 3'd1;
        frame3[6][16] = 3'd3;
        frame3[6][17] = 3'd3;
        frame3[6][18] = 3'd1;
        frame3[6][19] = 3'd1;
        frame3[6][20] = 3'd0;
        frame3[6][21] = 3'd0;
        frame3[6][22] = 3'd0;
        frame3[6][23] = 3'd0;
        frame3[6][24] = 3'd0;
        
        frame3[7][0] = 3'd0;
        frame3[7][1] = 3'd0;
        frame3[7][2] = 3'd0;
        frame3[7][3] = 3'd0;
        frame3[7][4] = 3'd0;
        frame3[7][5] = 3'd0;
        frame3[7][6] = 3'd0;
        frame3[7][7] = 3'd0;
        frame3[7][8] = 3'd0;
        frame3[7][9] = 3'd0;
        frame3[7][10] = 3'd0;
        frame3[7][11] = 3'd0;
        frame3[7][12] = 3'd0;
        frame3[7][13] = 3'd0;
        frame3[7][14] = 3'd0;
        frame3[7][15] = 3'd1;
        frame3[7][16] = 3'd2;
        frame3[7][17] = 3'd3;
        frame3[7][18] = 3'd1;
        frame3[7][19] = 3'd0;
        frame3[7][20] = 3'd0;
        frame3[7][21] = 3'd0;
        frame3[7][22] = 3'd0;
        frame3[7][23] = 3'd0;
        frame3[7][24] = 3'd0;
        
        frame3[8][0] = 3'd0;
        frame3[8][1] = 3'd0;
        frame3[8][2] = 3'd0;
        frame3[8][3] = 3'd0;
        frame3[8][4] = 3'd0;
        frame3[8][5] = 3'd0;
        frame3[8][6] = 3'd0;
        frame3[8][7] = 3'd0;
        frame3[8][8] = 3'd0;
        frame3[8][9] = 3'd0;
        frame3[8][10] = 3'd0;
        frame3[8][11] = 3'd0;
        frame3[8][12] = 3'd0;
        frame3[8][13] = 3'd0;
        frame3[8][14] = 3'd0;
        frame3[8][15] = 3'd1;
        frame3[8][16] = 3'd2;
        frame3[8][17] = 3'd2;
        frame3[8][18] = 3'd1;
        frame3[8][19] = 3'd0;
        frame3[8][20] = 3'd0;
        frame3[8][21] = 3'd0;
        frame3[8][22] = 3'd0;
        frame3[8][23] = 3'd0;
        frame3[8][24] = 3'd0;
        
        frame3[9][0] = 3'd0;
        frame3[9][1] = 3'd0;
        frame3[9][2] = 3'd0;
        frame3[9][3] = 3'd0;
        frame3[9][4] = 3'd0;
        frame3[9][5] = 3'd0;
        frame3[9][6] = 3'd0;
        frame3[9][7] = 3'd0;
        frame3[9][8] = 3'd0;
        frame3[9][9] = 3'd0;
        frame3[9][10] = 3'd0;
        frame3[9][11] = 3'd0;
        frame3[9][12] = 3'd0;
        frame3[9][13] = 3'd0;
        frame3[9][14] = 3'd0;
        frame3[9][15] = 3'd1;
        frame3[9][16] = 3'd2;
        frame3[9][17] = 3'd2;
        frame3[9][18] = 3'd1;
        frame3[9][19] = 3'd0;
        frame3[9][20] = 3'd0;
        frame3[9][21] = 3'd0;
        frame3[9][22] = 3'd0;
        frame3[9][23] = 3'd0;
        frame3[9][24] = 3'd0;
        
        frame3[10][0] = 3'd0;
        frame3[10][1] = 3'd0;
        frame3[10][2] = 3'd0;
        frame3[10][3] = 3'd0;
        frame3[10][4] = 3'd0;
        frame3[10][5] = 3'd0;
        frame3[10][6] = 3'd0;
        frame3[10][7] = 3'd0;
        frame3[10][8] = 3'd0;
        frame3[10][9] = 3'd0;
        frame3[10][10] = 3'd0;
        frame3[10][11] = 3'd0;
        frame3[10][12] = 3'd0;
        frame3[10][13] = 3'd0;
        frame3[10][14] = 3'd0;
        frame3[10][15] = 3'd1;
        frame3[10][16] = 3'd2;
        frame3[10][17] = 3'd2;
        frame3[10][18] = 3'd1;
        frame3[10][19] = 3'd0;
        frame3[10][20] = 3'd0;
        frame3[10][21] = 3'd0;
        frame3[10][22] = 3'd0;
        frame3[10][23] = 3'd0;
        frame3[10][24] = 3'd0;
        
        frame3[11][0] = 3'd0;
        frame3[11][1] = 3'd0;
        frame3[11][2] = 3'd0;
        frame3[11][3] = 3'd0;
        frame3[11][4] = 3'd0;
        frame3[11][5] = 3'd0;
        frame3[11][6] = 3'd0;
        frame3[11][7] = 3'd0;
        frame3[11][8] = 3'd0;
        frame3[11][9] = 3'd0;
        frame3[11][10] = 3'd0;
        frame3[11][11] = 3'd0;
        frame3[11][12] = 3'd0;
        frame3[11][13] = 3'd0;
        frame3[11][14] = 3'd1;
        frame3[11][15] = 3'd1;
        frame3[11][16] = 3'd2;
        frame3[11][17] = 3'd2;
        frame3[11][18] = 3'd1;
        frame3[11][19] = 3'd1;
        frame3[11][20] = 3'd0;
        frame3[11][21] = 3'd0;
        frame3[11][22] = 3'd0;
        frame3[11][23] = 3'd0;
        frame3[11][24] = 3'd0;
        
        frame3[12][0] = 3'd0;
        frame3[12][1] = 3'd1;
        frame3[12][2] = 3'd1;
        frame3[12][3] = 3'd0;
        frame3[12][4] = 3'd0;
        frame3[12][5] = 3'd0;
        frame3[12][6] = 3'd0;
        frame3[12][7] = 3'd0;
        frame3[12][8] = 3'd0;
        frame3[12][9] = 3'd1;
        frame3[12][10] = 3'd1;
        frame3[12][11] = 3'd1;
        frame3[12][12] = 3'd1;
        frame3[12][13] = 3'd1;
        frame3[12][14] = 3'd1;
        frame3[12][15] = 3'd2;
        frame3[12][16] = 3'd4;
        frame3[12][17] = 3'd4;
        frame3[12][18] = 3'd4;
        frame3[12][19] = 3'd1;
        frame3[12][20] = 3'd0;
        frame3[12][21] = 3'd0;
        frame3[12][22] = 3'd0;
        frame3[12][23] = 3'd0;
        frame3[12][24] = 3'd0;
        
        frame3[13][0] = 3'd0;
        frame3[13][1] = 3'd1;
        frame3[13][2] = 3'd5;
        frame3[13][3] = 3'd5;
        frame3[13][4] = 3'd1;
        frame3[13][5] = 3'd1;
        frame3[13][6] = 3'd1;
        frame3[13][7] = 3'd5;
        frame3[13][8] = 3'd5;
        frame3[13][9] = 3'd5;
        frame3[13][10] = 3'd5;
        frame3[13][11] = 3'd5;
        frame3[13][12] = 3'd5;
        frame3[13][13] = 3'd5;
        frame3[13][14] = 3'd5;
        frame3[13][15] = 3'd5;
        frame3[13][16] = 3'd5;
        frame3[13][17] = 3'd5;
        frame3[13][18] = 3'd4;
        frame3[13][19] = 3'd4;
        frame3[13][20] = 3'd1;
        frame3[13][21] = 3'd1;
        frame3[13][22] = 3'd0;
        frame3[13][23] = 3'd0;
        frame3[13][24] = 3'd0;
        
        frame3[14][0] = 3'd0;
        frame3[14][1] = 3'd1;
        frame3[14][2] = 3'd5;
        frame3[14][3] = 3'd5;
        frame3[14][4] = 3'd5;
        frame3[14][5] = 3'd5;
        frame3[14][6] = 3'd5;
        frame3[14][7] = 3'd5;
        frame3[14][8] = 3'd5;
        frame3[14][9] = 3'd5;
        frame3[14][10] = 3'd5;
        frame3[14][11] = 3'd5;
        frame3[14][12] = 3'd5;
        frame3[14][13] = 3'd2;
        frame3[14][14] = 3'd2;
        frame3[14][15] = 3'd5;
        frame3[14][16] = 3'd5;
        frame3[14][17] = 3'd5;
        frame3[14][18] = 3'd5;
        frame3[14][19] = 3'd4;
        frame3[14][20] = 3'd4;
        frame3[14][21] = 3'd1;
        frame3[14][22] = 3'd0;
        frame3[14][23] = 3'd0;
        frame3[14][24] = 3'd0;
        
        frame3[15][0] = 3'd0;
        frame3[15][1] = 3'd1;
        frame3[15][2] = 3'd5;
        frame3[15][3] = 3'd5;
        frame3[15][4] = 3'd5;
        frame3[15][5] = 3'd5;
        frame3[15][6] = 3'd5;
        frame3[15][7] = 3'd5;
        frame3[15][8] = 3'd5;
        frame3[15][9] = 3'd5;
        frame3[15][10] = 3'd5;
        frame3[15][11] = 3'd5;
        frame3[15][12] = 3'd5;
        frame3[15][13] = 3'd2;
        frame3[15][14] = 3'd1;
        frame3[15][15] = 3'd5;
        frame3[15][16] = 3'd5;
        frame3[15][17] = 3'd5;
        frame3[15][18] = 3'd5;
        frame3[15][19] = 3'd4;
        frame3[15][20] = 3'd4;
        frame3[15][21] = 3'd1;
        frame3[15][22] = 3'd0;
        frame3[15][23] = 3'd0;
        frame3[15][24] = 3'd0;
        
        frame3[16][0] = 3'd0;
        frame3[16][1] = 3'd0;
        frame3[16][2] = 3'd1;
        frame3[16][3] = 3'd1;
        frame3[16][4] = 3'd3;
        frame3[16][5] = 3'd2;
        frame3[16][6] = 3'd2;
        frame3[16][7] = 3'd2;
        frame3[16][8] = 3'd2;
        frame3[16][9] = 3'd2;
        frame3[16][10] = 3'd2;
        frame3[16][11] = 3'd2;
        frame3[16][12] = 3'd1;
        frame3[16][13] = 3'd5;
        frame3[16][14] = 3'd5;
        frame3[16][15] = 3'd5;
        frame3[16][16] = 3'd5;
        frame3[16][17] = 3'd5;
        frame3[16][18] = 3'd4;
        frame3[16][19] = 3'd4;
        frame3[16][20] = 3'd4;
        frame3[16][21] = 3'd1;
        frame3[16][22] = 3'd0;
        frame3[16][23] = 3'd0;
        frame3[16][24] = 3'd0;
        
        frame3[17][0] = 3'd0;
        frame3[17][1] = 3'd0;
        frame3[17][2] = 3'd0;
        frame3[17][3] = 3'd1;
        frame3[17][4] = 3'd1;
        frame3[17][5] = 3'd1;
        frame3[17][6] = 3'd1;
        frame3[17][7] = 3'd1;
        frame3[17][8] = 3'd1;
        frame3[17][9] = 3'd1;
        frame3[17][10] = 3'd1;
        frame3[17][11] = 3'd1;
        frame3[17][12] = 3'd5;
        frame3[17][13] = 3'd5;
        frame3[17][14] = 3'd5;
        frame3[17][15] = 3'd5;
        frame3[17][16] = 3'd5;
        frame3[17][17] = 3'd4;
        frame3[17][18] = 3'd4;
        frame3[17][19] = 3'd4;
        frame3[17][20] = 3'd1;
        frame3[17][21] = 3'd1;
        frame3[17][22] = 3'd0;
        frame3[17][23] = 3'd0;
        frame3[17][24] = 3'd0;
        
        frame3[18][0] = 3'd0;
        frame3[18][1] = 3'd0;
        frame3[18][2] = 3'd0;
        frame3[18][3] = 3'd0;
        frame3[18][4] = 3'd1;
        frame3[18][5] = 3'd3;
        frame3[18][6] = 3'd3;
        frame3[18][7] = 3'd3;
        frame3[18][8] = 3'd3;
        frame3[18][9] = 3'd3;
        frame3[18][10] = 3'd3;
        frame3[18][11] = 3'd3;
        frame3[18][12] = 3'd5;
        frame3[18][13] = 3'd5;
        frame3[18][14] = 3'd5;
        frame3[18][15] = 3'd5;
        frame3[18][16] = 3'd4;
        frame3[18][17] = 3'd4;
        frame3[18][18] = 3'd4;
        frame3[18][19] = 3'd1;
        frame3[18][20] = 3'd0;
        frame3[18][21] = 3'd0;
        frame3[18][22] = 3'd0;
        frame3[18][23] = 3'd0;
        frame3[18][24] = 3'd0;
        
        frame3[19][0] = 3'd0;
        frame3[19][1] = 3'd0;
        frame3[19][2] = 3'd0;
        frame3[19][3] = 3'd0;
        frame3[19][4] = 3'd0;
        frame3[19][5] = 3'd1;
        frame3[19][6] = 3'd4;
        frame3[19][7] = 3'd4;
        frame3[19][8] = 3'd3;
        frame3[19][9] = 3'd3;
        frame3[19][10] = 3'd3;
        frame3[19][11] = 3'd4;
        frame3[19][12] = 3'd4;
        frame3[19][13] = 3'd4;
        frame3[19][14] = 3'd4;
        frame3[19][15] = 3'd4;
        frame3[19][16] = 3'd4;
        frame3[19][17] = 3'd4;
        frame3[19][18] = 3'd1;
        frame3[19][19] = 3'd1;
        frame3[19][20] = 3'd0;
        frame3[19][21] = 3'd0;
        frame3[19][22] = 3'd0;
        frame3[19][23] = 3'd0;
        frame3[19][24] = 3'd0;
        
        frame3[20][0] = 3'd0;
        frame3[20][1] = 3'd0;
        frame3[20][2] = 3'd0;
        frame3[20][3] = 3'd0;
        frame3[20][4] = 3'd0;
        frame3[20][5] = 3'd0;
        frame3[20][6] = 3'd0;
        frame3[20][7] = 3'd1;
        frame3[20][8] = 3'd1;
        frame3[20][9] = 3'd1;
        frame3[20][10] = 3'd1;
        frame3[20][11] = 3'd1;
        frame3[20][12] = 3'd5;
        frame3[20][13] = 3'd5;
        frame3[20][14] = 3'd1;
        frame3[20][15] = 3'd1;
        frame3[20][16] = 3'd1;
        frame3[20][17] = 3'd0;
        frame3[20][18] = 3'd0;
        frame3[20][19] = 3'd0;
        frame3[20][20] = 3'd0;
        frame3[20][21] = 3'd0;
        frame3[20][22] = 3'd0;
        frame3[20][23] = 3'd0;
        frame3[20][24] = 3'd0;
        
        frame3[21][0] = 3'd0;
        frame3[21][1] = 3'd0;
        frame3[21][2] = 3'd0;
        frame3[21][3] = 3'd0;
        frame3[21][4] = 3'd0;
        frame3[21][5] = 3'd0;
        frame3[21][6] = 3'd0;
        frame3[21][7] = 3'd0;
        frame3[21][8] = 3'd0;
        frame3[21][9] = 3'd1;
        frame3[21][10] = 3'd0;
        frame3[21][11] = 3'd1;
        frame3[21][12] = 3'd1;
        frame3[21][13] = 3'd1;
        frame3[21][14] = 3'd1;
        frame3[21][15] = 3'd0;
        frame3[21][16] = 3'd0;
        frame3[21][17] = 3'd0;
        frame3[21][18] = 3'd0;
        frame3[21][19] = 3'd0;
        frame3[21][20] = 3'd0;
        frame3[21][21] = 3'd0;
        frame3[21][22] = 3'd0;
        frame3[21][23] = 3'd0;
        frame3[21][24] = 3'd0;
        
        frame3[22][0] = 3'd0;
        frame3[22][1] = 3'd0;
        frame3[22][2] = 3'd0;
        frame3[22][3] = 3'd0;
        frame3[22][4] = 3'd0;
        frame3[22][5] = 3'd0;
        frame3[22][6] = 3'd0;
        frame3[22][7] = 3'd0;
        frame3[22][8] = 3'd0;
        frame3[22][9] = 3'd1;
        frame3[22][10] = 3'd0;
        frame3[22][11] = 3'd0;
        frame3[22][12] = 3'd0;
        frame3[22][13] = 3'd1;
        frame3[22][14] = 3'd0;
        frame3[22][15] = 3'd0;
        frame3[22][16] = 3'd0;
        frame3[22][17] = 3'd0;
        frame3[22][18] = 3'd0;
        frame3[22][19] = 3'd0;
        frame3[22][20] = 3'd0;
        frame3[22][21] = 3'd0;
        frame3[22][22] = 3'd0;
        frame3[22][23] = 3'd0;
        frame3[22][24] = 3'd0;
        
        frame3[23][0] = 3'd0;
        frame3[23][1] = 3'd0;
        frame3[23][2] = 3'd0;
        frame3[23][3] = 3'd0;
        frame3[23][4] = 3'd0;
        frame3[23][5] = 3'd0;
        frame3[23][6] = 3'd0;
        frame3[23][7] = 3'd0;
        frame3[23][8] = 3'd0;
        frame3[23][9] = 3'd1;
        frame3[23][10] = 3'd1;
        frame3[23][11] = 3'd0;
        frame3[23][12] = 3'd0;
        frame3[23][13] = 3'd1;
        frame3[23][14] = 3'd1;
        frame3[23][15] = 3'd0;
        frame3[23][16] = 3'd0;
        frame3[23][17] = 3'd0;
        frame3[23][18] = 3'd0;
        frame3[23][19] = 3'd0;
        frame3[23][20] = 3'd0;
        frame3[23][21] = 3'd0;
        frame3[23][22] = 3'd0;
        frame3[23][23] = 3'd0;
        frame3[23][24] = 3'd0;
        
        frame3[24][0] = 3'd0;
        frame3[24][1] = 3'd0;
        frame3[24][2] = 3'd0;
        frame3[24][3] = 3'd0;
        frame3[24][4] = 3'd0;
        frame3[24][5] = 3'd0;
        frame3[24][6] = 3'd0;
        frame3[24][7] = 3'd0;
        frame3[24][8] = 3'd0;
        frame3[24][9] = 3'd1;
        frame3[24][10] = 3'd1;
        frame3[24][11] = 3'd1;
        frame3[24][12] = 3'd0;
        frame3[24][13] = 3'd1;
        frame3[24][14] = 3'd1;
        frame3[24][15] = 3'd1;
        frame3[24][16] = 3'd0;
        frame3[24][17] = 3'd0;
        frame3[24][18] = 3'd0;
        frame3[24][19] = 3'd0;
        frame3[24][20] = 3'd0;
        frame3[24][21] = 3'd0;
        frame3[24][22] = 3'd0;
        frame3[24][23] = 3'd0;
        frame3[24][24] = 3'd0;
    end