reg [2:0] frame2 [0:24][0:24] = '{
    '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,2,2,2,2,2,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,2,2,2,2,2,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,4,2,2,2,4,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,0,1,1,2,1,1,0,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,0,0,1,2,1,0,0,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,0,0,1,2,1,0,0,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,0,0,1,2,1,0,0,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,0,0,1,2,1,0,0,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,1,1,2,1,1,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,5,5,5,5,5,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,1,5,5,5,5,5,5,5,1,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,1,1,5,5,5,5,5,5,5,5,5,1,1,0,0,0,0,0,0},
    '{0,0,0,0,0,1,1,2,5,5,5,5,5,5,5,5,5,2,1,1,0,0,0,0,0},
    '{0,0,0,0,0,1,2,2,5,5,5,5,5,5,5,5,5,2,2,1,0,0,0,0,0},
    '{0,0,0,0,0,1,1,1,1,2,5,5,5,5,5,2,1,1,1,1,0,0,0,0,0},
    '{0,0,0,0,0,0,1,3,4,1,2,2,5,2,2,1,4,3,1,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,1,3,1,1,1,2,1,1,1,3,1,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,1,4,4,1,1,1,4,4,1,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,1,3,4,3,1,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,0,1,1,1,0,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0},
    '{0,0,0,0,0,0,0,0,1,1,0,1,0,1,0,1,1,0,0,0,0,0,0,0,0}
};
