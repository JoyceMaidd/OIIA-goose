reg [2:0] frame2 [0:1][0:1];

initial begin
    frame2[0][0] = 3'h0;
    frame2[0][1] = 3'h0;
    // frame2[0][2] = 3'h0;
    // frame2[0][3] = 3'h0;
    // frame2[0][4] = 3'h0;
    // frame2[0][5] = 3'h0;
    // frame2[0][6] = 3'h0;
    // frame2[0][7] = 3'h0;
    // frame2[0][8] = 3'h0;
    // frame2[0][9] = 3'h0;
    // frame2[0][10] = 3'h0;
    // frame2[0][11] = 3'h0;
    // frame2[0][12] = 3'h0;
    // frame2[0][13] = 3'h0;
    // frame2[0][14] = 3'h0;
    // frame2[0][15] = 3'h0;
    // frame2[0][16] = 3'h0;
    // frame2[0][17] = 3'h0;
    // frame2[0][18] = 3'h0;
    // frame2[0][19] = 3'h0;
    // frame2[0][20] = 3'h0;
    // frame2[0][21] = 3'h0;
    // frame2[0][22] = 3'h0;
    // frame2[0][23] = 3'h0;
    // frame2[0][24] = 3'h0;
    // frame2[0][25] = 3'h0;
    // frame2[0][26] = 3'h0;
    // frame2[0][27] = 3'h0;
    // frame2[0][28] = 3'h0;
    // frame2[0][29] = 3'h0;
    // frame2[0][30] = 3'h0;
    // frame2[0][31] = 3'h0;
    frame2[1][0] = 3'h0;
    frame2[1][1] = 3'h0;
    // frame2[1][2] = 3'h0;
    // frame2[1][3] = 3'h0;
    // frame2[1][4] = 3'h0;
    // frame2[1][5] = 3'h0;
    // frame2[1][6] = 3'h0;
    // frame2[1][7] = 3'h0;
    // frame2[1][8] = 3'h0;
    // frame2[1][9] = 3'h0;
    // frame2[1][10] = 3'h0;
    // frame2[1][11] = 3'h0;
    // frame2[1][12] = 3'h0;
    // frame2[1][13] = 3'h1;
    // frame2[1][14] = 3'h1;
    // frame2[1][15] = 3'h1;
    // frame2[1][16] = 3'h1;
    // frame2[1][17] = 3'h1;
    // frame2[1][18] = 3'h1;
    // frame2[1][19] = 3'h0;
    // frame2[1][20] = 3'h0;
    // frame2[1][21] = 3'h0;
    // frame2[1][22] = 3'h0;
    // frame2[1][23] = 3'h0;
    // frame2[1][24] = 3'h0;
    // frame2[1][25] = 3'h0;
    // frame2[1][26] = 3'h0;
    // frame2[1][27] = 3'h0;
    // frame2[1][28] = 3'h0;
    // frame2[1][29] = 3'h0;
    // frame2[1][30] = 3'h0;
    // frame2[1][31] = 3'h0;
    // frame2[2][0] = 3'h0;
    // frame2[2][1] = 3'h0;
    // frame2[2][2] = 3'h0;
    // frame2[2][3] = 3'h0;
    // frame2[2][4] = 3'h0;
    // frame2[2][5] = 3'h0;
    // frame2[2][6] = 3'h0;
    // frame2[2][7] = 3'h0;
    // frame2[2][8] = 3'h0;
    // frame2[2][9] = 3'h0;
    // frame2[2][10] = 3'h0;
    // frame2[2][11] = 3'h0;
    // frame2[2][12] = 3'h1;
    // frame2[2][13] = 3'h1;
    // frame2[2][14] = 3'h2;
    // frame2[2][15] = 3'h2;
    // frame2[2][16] = 3'h2;
    // frame2[2][17] = 3'h2;
    // frame2[2][18] = 3'h1;
    // frame2[2][19] = 3'h1;
    // frame2[2][20] = 3'h0;
    // frame2[2][21] = 3'h0;
    // frame2[2][22] = 3'h0;
    // frame2[2][23] = 3'h0;
    // frame2[2][24] = 3'h0;
    // frame2[2][25] = 3'h0;
    // frame2[2][26] = 3'h0;
    // frame2[2][27] = 3'h0;
    // frame2[2][28] = 3'h0;
    // frame2[2][29] = 3'h0;
    // frame2[2][30] = 3'h0;
    // frame2[2][31] = 3'h0;
    // frame2[3][0] = 3'h0;
    // frame2[3][1] = 3'h0;
    // frame2[3][2] = 3'h0;
    // frame2[3][3] = 3'h0;
    // frame2[3][4] = 3'h0;
    // frame2[3][5] = 3'h0;
    // frame2[3][6] = 3'h0;
    // frame2[3][7] = 3'h0;
    // frame2[3][8] = 3'h0;
    // frame2[3][9] = 3'h0;
    // frame2[3][10] = 3'h0;
    // frame2[3][11] = 3'h0;
    // frame2[3][12] = 3'h1;
    // frame2[3][13] = 3'h2;
    // frame2[3][14] = 3'h2;
    // frame2[3][15] = 3'h2;
    // frame2[3][16] = 3'h2;
    // frame2[3][17] = 3'h2;
    // frame2[3][18] = 3'h2;
    // frame2[3][19] = 3'h1;
    // frame2[3][20] = 3'h0;
    // frame2[3][21] = 3'h0;
    // frame2[3][22] = 3'h0;
    // frame2[3][23] = 3'h0;
    // frame2[3][24] = 3'h0;
    // frame2[3][25] = 3'h0;
    // frame2[3][26] = 3'h0;
    // frame2[3][27] = 3'h0;
    // frame2[3][28] = 3'h0;
    // frame2[3][29] = 3'h0;
    // frame2[3][30] = 3'h0;
    // frame2[3][31] = 3'h0;
    // frame2[4][0] = 3'h0;
    // frame2[4][1] = 3'h0;
    // frame2[4][2] = 3'h0;
    // frame2[4][3] = 3'h0;
    // frame2[4][4] = 3'h0;
    // frame2[4][5] = 3'h0;
    // frame2[4][6] = 3'h0;
    // frame2[4][7] = 3'h0;
    // frame2[4][8] = 3'h0;
    // frame2[4][9] = 3'h0;
    // frame2[4][10] = 3'h0;
    // frame2[4][11] = 3'h0;
    // frame2[4][12] = 3'h1;
    // frame2[4][13] = 3'h2;
    // frame2[4][14] = 3'h2;
    // frame2[4][15] = 3'h2;
    // frame2[4][16] = 3'h2;
    // frame2[4][17] = 3'h2;
    // frame2[4][18] = 3'h2;
    // frame2[4][19] = 3'h1;
    // frame2[4][20] = 3'h0;
    // frame2[4][21] = 3'h0;
    // frame2[4][22] = 3'h0;
    // frame2[4][23] = 3'h0;
    // frame2[4][24] = 3'h0;
    // frame2[4][25] = 3'h0;
    // frame2[4][26] = 3'h0;
    // frame2[4][27] = 3'h0;
    // frame2[4][28] = 3'h0;
    // frame2[4][29] = 3'h0;
    // frame2[4][30] = 3'h0;
    // frame2[4][31] = 3'h0;
    // frame2[5][0] = 3'h0;
    // frame2[5][1] = 3'h0;
    // frame2[5][2] = 3'h0;
    // frame2[5][3] = 3'h0;
    // frame2[5][4] = 3'h0;
    // frame2[5][5] = 3'h0;
    // frame2[5][6] = 3'h0;
    // frame2[5][7] = 3'h0;
    // frame2[5][8] = 3'h0;
    // frame2[5][9] = 3'h0;
    // frame2[5][10] = 3'h0;
    // frame2[5][11] = 3'h0;
    // frame2[5][12] = 3'h1;
    // frame2[5][13] = 3'h4;
    // frame2[5][14] = 3'h2;
    // frame2[5][15] = 3'h2;
    // frame2[5][16] = 3'h2;
    // frame2[5][17] = 3'h2;
    // frame2[5][18] = 3'h4;
    // frame2[5][19] = 3'h1;
    // frame2[5][20] = 3'h0;
    // frame2[5][21] = 3'h0;
    // frame2[5][22] = 3'h0;
    // frame2[5][23] = 3'h0;
    // frame2[5][24] = 3'h0;
    // frame2[5][25] = 3'h0;
    // frame2[5][26] = 3'h0;
    // frame2[5][27] = 3'h0;
    // frame2[5][28] = 3'h0;
    // frame2[5][29] = 3'h0;
    // frame2[5][30] = 3'h0;
    // frame2[5][31] = 3'h0;
    // frame2[6][0] = 3'h0;
    // frame2[6][1] = 3'h0;
    // frame2[6][2] = 3'h0;
    // frame2[6][3] = 3'h0;
    // frame2[6][4] = 3'h0;
    // frame2[6][5] = 3'h0;
    // frame2[6][6] = 3'h0;
    // frame2[6][7] = 3'h0;
    // frame2[6][8] = 3'h0;
    // frame2[6][9] = 3'h0;
    // frame2[6][10] = 3'h0;
    // frame2[6][11] = 3'h0;
    // frame2[6][12] = 3'h1;
    // frame2[6][13] = 3'h1;
    // frame2[6][14] = 3'h4;
    // frame2[6][15] = 3'h2;
    // frame2[6][16] = 3'h2;
    // frame2[6][17] = 3'h4;
    // frame2[6][18] = 3'h1;
    // frame2[6][19] = 3'h1;
    // frame2[6][20] = 3'h0;
    // frame2[6][21] = 3'h0;
    // frame2[6][22] = 3'h0;
    // frame2[6][23] = 3'h0;
    // frame2[6][24] = 3'h0;
    // frame2[6][25] = 3'h0;
    // frame2[6][26] = 3'h0;
    // frame2[6][27] = 3'h0;
    // frame2[6][28] = 3'h0;
    // frame2[6][29] = 3'h0;
    // frame2[6][30] = 3'h0;
    // frame2[6][31] = 3'h0;
    // frame2[7][0] = 3'h0;
    // frame2[7][1] = 3'h0;
    // frame2[7][2] = 3'h0;
    // frame2[7][3] = 3'h0;
    // frame2[7][4] = 3'h0;
    // frame2[7][5] = 3'h0;
    // frame2[7][6] = 3'h0;
    // frame2[7][7] = 3'h0;
    // frame2[7][8] = 3'h0;
    // frame2[7][9] = 3'h0;
    // frame2[7][10] = 3'h0;
    // frame2[7][11] = 3'h0;
    // frame2[7][12] = 3'h0;
    // frame2[7][13] = 3'h1;
    // frame2[7][14] = 3'h1;
    // frame2[7][15] = 3'h2;
    // frame2[7][16] = 3'h2;
    // frame2[7][17] = 3'h1;
    // frame2[7][18] = 3'h1;
    // frame2[7][19] = 3'h0;
    // frame2[7][20] = 3'h0;
    // frame2[7][21] = 3'h0;
    // frame2[7][22] = 3'h0;
    // frame2[7][23] = 3'h0;
    // frame2[7][24] = 3'h0;
    // frame2[7][25] = 3'h0;
    // frame2[7][26] = 3'h0;
    // frame2[7][27] = 3'h0;
    // frame2[7][28] = 3'h0;
    // frame2[7][29] = 3'h0;
    // frame2[7][30] = 3'h0;
    // frame2[7][31] = 3'h0;
    // frame2[8][0] = 3'h0;
    // frame2[8][1] = 3'h0;
    // frame2[8][2] = 3'h0;
    // frame2[8][3] = 3'h0;
    // frame2[8][4] = 3'h0;
    // frame2[8][5] = 3'h0;
    // frame2[8][6] = 3'h0;
    // frame2[8][7] = 3'h0;
    // frame2[8][8] = 3'h0;
    // frame2[8][9] = 3'h0;
    // frame2[8][10] = 3'h0;
    // frame2[8][11] = 3'h0;
    // frame2[8][12] = 3'h0;
    // frame2[8][13] = 3'h0;
    // frame2[8][14] = 3'h1;
    // frame2[8][15] = 3'h2;
    // frame2[8][16] = 3'h2;
    // frame2[8][17] = 3'h1;
    // frame2[8][18] = 3'h0;
    // frame2[8][19] = 3'h0;
    // frame2[8][20] = 3'h0;
    // frame2[8][21] = 3'h0;
    // frame2[8][22] = 3'h0;
    // frame2[8][23] = 3'h0;
    // frame2[8][24] = 3'h0;
    // frame2[8][25] = 3'h0;
    // frame2[8][26] = 3'h0;
    // frame2[8][27] = 3'h0;
    // frame2[8][28] = 3'h0;
    // frame2[8][29] = 3'h0;
    // frame2[8][30] = 3'h0;
    // frame2[8][31] = 3'h0;
    // frame2[9][0] = 3'h0;
    // frame2[9][1] = 3'h0;
    // frame2[9][2] = 3'h0;
    // frame2[9][3] = 3'h0;
    // frame2[9][4] = 3'h0;
    // frame2[9][5] = 3'h0;
    // frame2[9][6] = 3'h0;
    // frame2[9][7] = 3'h0;
    // frame2[9][8] = 3'h0;
    // frame2[9][9] = 3'h0;
    // frame2[9][10] = 3'h0;
    // frame2[9][11] = 3'h0;
    // frame2[9][12] = 3'h0;
    // frame2[9][13] = 3'h0;
    // frame2[9][14] = 3'h1;
    // frame2[9][15] = 3'h2;
    // frame2[9][16] = 3'h2;
    // frame2[9][17] = 3'h1;
    // frame2[9][18] = 3'h0;
    // frame2[9][19] = 3'h0;
    // frame2[9][20] = 3'h0;
    // frame2[9][21] = 3'h0;
    // frame2[9][22] = 3'h0;
    // frame2[9][23] = 3'h0;
    // frame2[9][24] = 3'h0;
    // frame2[9][25] = 3'h0;
    // frame2[9][26] = 3'h0;
    // frame2[9][27] = 3'h0;
    // frame2[9][28] = 3'h0;
    // frame2[9][29] = 3'h0;
    // frame2[9][30] = 3'h0;
    // frame2[9][31] = 3'h0;
    // frame2[10][0] = 3'h0;
    // frame2[10][1] = 3'h0;
    // frame2[10][2] = 3'h0;
    // frame2[10][3] = 3'h0;
    // frame2[10][4] = 3'h0;
    // frame2[10][5] = 3'h0;
    // frame2[10][6] = 3'h0;
    // frame2[10][7] = 3'h0;
    // frame2[10][8] = 3'h0;
    // frame2[10][9] = 3'h0;
    // frame2[10][10] = 3'h0;
    // frame2[10][11] = 3'h0;
    // frame2[10][12] = 3'h0;
    // frame2[10][13] = 3'h0;
    // frame2[10][14] = 3'h1;
    // frame2[10][15] = 3'h2;
    // frame2[10][16] = 3'h2;
    // frame2[10][17] = 3'h1;
    // frame2[10][18] = 3'h0;
    // frame2[10][19] = 3'h0;
    // frame2[10][20] = 3'h0;
    // frame2[10][21] = 3'h0;
    // frame2[10][22] = 3'h0;
    // frame2[10][23] = 3'h0;
    // frame2[10][24] = 3'h0;
    // frame2[10][25] = 3'h0;
    // frame2[10][26] = 3'h0;
    // frame2[10][27] = 3'h0;
    // frame2[10][28] = 3'h0;
    // frame2[10][29] = 3'h0;
    // frame2[10][30] = 3'h0;
    // frame2[10][31] = 3'h0;
    // frame2[11][0] = 3'h0;
    // frame2[11][1] = 3'h0;
    // frame2[11][2] = 3'h0;
    // frame2[11][3] = 3'h0;
    // frame2[11][4] = 3'h0;
    // frame2[11][5] = 3'h0;
    // frame2[11][6] = 3'h0;
    // frame2[11][7] = 3'h0;
    // frame2[11][8] = 3'h0;
    // frame2[11][9] = 3'h0;
    // frame2[11][10] = 3'h0;
    // frame2[11][11] = 3'h0;
    // frame2[11][12] = 3'h0;
    // frame2[11][13] = 3'h0;
    // frame2[11][14] = 3'h1;
    // frame2[11][15] = 3'h2;
    // frame2[11][16] = 3'h2;
    // frame2[11][17] = 3'h1;
    // frame2[11][18] = 3'h0;
    // frame2[11][19] = 3'h0;
    // frame2[11][20] = 3'h0;
    // frame2[11][21] = 3'h0;
    // frame2[11][22] = 3'h0;
    // frame2[11][23] = 3'h0;
    // frame2[11][24] = 3'h0;
    // frame2[11][25] = 3'h0;
    // frame2[11][26] = 3'h0;
    // frame2[11][27] = 3'h0;
    // frame2[11][28] = 3'h0;
    // frame2[11][29] = 3'h0;
    // frame2[11][30] = 3'h0;
    // frame2[11][31] = 3'h0;
    // frame2[12][0] = 3'h0;
    // frame2[12][1] = 3'h0;
    // frame2[12][2] = 3'h0;
    // frame2[12][3] = 3'h0;
    // frame2[12][4] = 3'h0;
    // frame2[12][5] = 3'h0;
    // frame2[12][6] = 3'h0;
    // frame2[12][7] = 3'h0;
    // frame2[12][8] = 3'h0;
    // frame2[12][9] = 3'h0;
    // frame2[12][10] = 3'h0;
    // frame2[12][11] = 3'h0;
    // frame2[12][12] = 3'h0;
    // frame2[12][13] = 3'h0;
    // frame2[12][14] = 3'h1;
    // frame2[12][15] = 3'h2;
    // frame2[12][16] = 3'h2;
    // frame2[12][17] = 3'h1;
    // frame2[12][18] = 3'h0;
    // frame2[12][19] = 3'h0;
    // frame2[12][20] = 3'h0;
    // frame2[12][21] = 3'h0;
    // frame2[12][22] = 3'h0;
    // frame2[12][23] = 3'h0;
    // frame2[12][24] = 3'h0;
    // frame2[12][25] = 3'h0;
    // frame2[12][26] = 3'h0;
    // frame2[12][27] = 3'h0;
    // frame2[12][28] = 3'h0;
    // frame2[12][29] = 3'h0;
    // frame2[12][30] = 3'h0;
    // frame2[12][31] = 3'h0;
    // frame2[13][0] = 3'h0;
    // frame2[13][1] = 3'h0;
    // frame2[13][2] = 3'h0;
    // frame2[13][3] = 3'h0;
    // frame2[13][4] = 3'h0;
    // frame2[13][5] = 3'h0;
    // frame2[13][6] = 3'h0;
    // frame2[13][7] = 3'h0;
    // frame2[13][8] = 3'h0;
    // frame2[13][9] = 3'h0;
    // frame2[13][10] = 3'h0;
    // frame2[13][11] = 3'h0;
    // frame2[13][12] = 3'h1;
    // frame2[13][13] = 3'h1;
    // frame2[13][14] = 3'h1;
    // frame2[13][15] = 3'h2;
    // frame2[13][16] = 3'h2;
    // frame2[13][17] = 3'h1;
    // frame2[13][18] = 3'h1;
    // frame2[13][19] = 3'h1;
    // frame2[13][20] = 3'h0;
    // frame2[13][21] = 3'h0;
    // frame2[13][22] = 3'h0;
    // frame2[13][23] = 3'h0;
    // frame2[13][24] = 3'h0;
    // frame2[13][25] = 3'h0;
    // frame2[13][26] = 3'h0;
    // frame2[13][27] = 3'h0;
    // frame2[13][28] = 3'h0;
    // frame2[13][29] = 3'h0;
    // frame2[13][30] = 3'h0;
    // frame2[13][31] = 3'h0;
    // frame2[14][0] = 3'h0;
    // frame2[14][1] = 3'h0;
    // frame2[14][2] = 3'h0;
    // frame2[14][3] = 3'h0;
    // frame2[14][4] = 3'h0;
    // frame2[14][5] = 3'h0;
    // frame2[14][6] = 3'h0;
    // frame2[14][7] = 3'h0;
    // frame2[14][8] = 3'h0;
    // frame2[14][9] = 3'h0;
    // frame2[14][10] = 3'h0;
    // frame2[14][11] = 3'h1;
    // frame2[14][12] = 3'h1;
    // frame2[14][13] = 3'h5;
    // frame2[14][14] = 3'h5;
    // frame2[14][15] = 3'h5;
    // frame2[14][16] = 3'h5;
    // frame2[14][17] = 3'h5;
    // frame2[14][18] = 3'h5;
    // frame2[14][19] = 3'h1;
    // frame2[14][20] = 3'h1;
    // frame2[14][21] = 3'h0;
    // frame2[14][22] = 3'h0;
    // frame2[14][23] = 3'h0;
    // frame2[14][24] = 3'h0;
    // frame2[14][25] = 3'h0;
    // frame2[14][26] = 3'h0;
    // frame2[14][27] = 3'h0;
    // frame2[14][28] = 3'h0;
    // frame2[14][29] = 3'h0;
    // frame2[14][30] = 3'h0;
    // frame2[14][31] = 3'h0;
    // frame2[15][0] = 3'h0;
    // frame2[15][1] = 3'h0;
    // frame2[15][2] = 3'h0;
    // frame2[15][3] = 3'h0;
    // frame2[15][4] = 3'h0;
    // frame2[15][5] = 3'h0;
    // frame2[15][6] = 3'h0;
    // frame2[15][7] = 3'h0;
    // frame2[15][8] = 3'h0;
    // frame2[15][9] = 3'h0;
    // frame2[15][10] = 3'h1;
    // frame2[15][11] = 3'h1;
    // frame2[15][12] = 3'h5;
    // frame2[15][13] = 3'h5;
    // frame2[15][14] = 3'h5;
    // frame2[15][15] = 3'h5;
    // frame2[15][16] = 3'h5;
    // frame2[15][17] = 3'h5;
    // frame2[15][18] = 3'h5;
    // frame2[15][19] = 3'h5;
    // frame2[15][20] = 3'h1;
    // frame2[15][21] = 3'h1;
    // frame2[15][22] = 3'h0;
    // frame2[15][23] = 3'h0;
    // frame2[15][24] = 3'h0;
    // frame2[15][25] = 3'h0;
    // frame2[15][26] = 3'h0;
    // frame2[15][27] = 3'h0;
    // frame2[15][28] = 3'h0;
    // frame2[15][29] = 3'h0;
    // frame2[15][30] = 3'h0;
    // frame2[15][31] = 3'h0;
    // frame2[16][0] = 3'h0;
    // frame2[16][1] = 3'h0;
    // frame2[16][2] = 3'h0;
    // frame2[16][3] = 3'h0;
    // frame2[16][4] = 3'h0;
    // frame2[16][5] = 3'h0;
    // frame2[16][6] = 3'h0;
    // frame2[16][7] = 3'h0;
    // frame2[16][8] = 3'h0;
    // frame2[16][9] = 3'h1;
    // frame2[16][10] = 3'h1;
    // frame2[16][11] = 3'h5;
    // frame2[16][12] = 3'h5;
    // frame2[16][13] = 3'h5;
    // frame2[16][14] = 3'h5;
    // frame2[16][15] = 3'h5;
    // frame2[16][16] = 3'h5;
    // frame2[16][17] = 3'h5;
    // frame2[16][18] = 3'h5;
    // frame2[16][19] = 3'h5;
    // frame2[16][20] = 3'h5;
    // frame2[16][21] = 3'h1;
    // frame2[16][22] = 3'h1;
    // frame2[16][23] = 3'h0;
    // frame2[16][24] = 3'h0;
    // frame2[16][25] = 3'h0;
    // frame2[16][26] = 3'h0;
    // frame2[16][27] = 3'h0;
    // frame2[16][28] = 3'h0;
    // frame2[16][29] = 3'h0;
    // frame2[16][30] = 3'h0;
    // frame2[16][31] = 3'h0;
    // frame2[17][0] = 3'h0;
    // frame2[17][1] = 3'h0;
    // frame2[17][2] = 3'h0;
    // frame2[17][3] = 3'h0;
    // frame2[17][4] = 3'h0;
    // frame2[17][5] = 3'h0;
    // frame2[17][6] = 3'h0;
    // frame2[17][7] = 3'h0;
    // frame2[17][8] = 3'h1;
    // frame2[17][9] = 3'h1;
    // frame2[17][10] = 3'h5;
    // frame2[17][11] = 3'h5;
    // frame2[17][12] = 3'h5;
    // frame2[17][13] = 3'h5;
    // frame2[17][14] = 3'h5;
    // frame2[17][15] = 3'h5;
    // frame2[17][16] = 3'h5;
    // frame2[17][17] = 3'h5;
    // frame2[17][18] = 3'h5;
    // frame2[17][19] = 3'h5;
    // frame2[17][20] = 3'h5;
    // frame2[17][21] = 3'h5;
    // frame2[17][22] = 3'h1;
    // frame2[17][23] = 3'h1;
    // frame2[17][24] = 3'h0;
    // frame2[17][25] = 3'h0;
    // frame2[17][26] = 3'h0;
    // frame2[17][27] = 3'h0;
    // frame2[17][28] = 3'h0;
    // frame2[17][29] = 3'h0;
    // frame2[17][30] = 3'h0;
    // frame2[17][31] = 3'h0;
    // frame2[18][0] = 3'h0;
    // frame2[18][1] = 3'h0;
    // frame2[18][2] = 3'h0;
    // frame2[18][3] = 3'h0;
    // frame2[18][4] = 3'h0;
    // frame2[18][5] = 3'h0;
    // frame2[18][6] = 3'h0;
    // frame2[18][7] = 3'h1;
    // frame2[18][8] = 3'h1;
    // frame2[18][9] = 3'h2;
    // frame2[18][10] = 3'h5;
    // frame2[18][11] = 3'h5;
    // frame2[18][12] = 3'h5;
    // frame2[18][13] = 3'h5;
    // frame2[18][14] = 3'h5;
    // frame2[18][15] = 3'h5;
    // frame2[18][16] = 3'h5;
    // frame2[18][17] = 3'h5;
    // frame2[18][18] = 3'h5;
    // frame2[18][19] = 3'h5;
    // frame2[18][20] = 3'h5;
    // frame2[18][21] = 3'h5;
    // frame2[18][22] = 3'h2;
    // frame2[18][23] = 3'h1;
    // frame2[18][24] = 3'h1;
    // frame2[18][25] = 3'h0;
    // frame2[18][26] = 3'h0;
    // frame2[18][27] = 3'h0;
    // frame2[18][28] = 3'h0;
    // frame2[18][29] = 3'h0;
    // frame2[18][30] = 3'h0;
    // frame2[18][31] = 3'h0;
    // frame2[19][0] = 3'h0;
    // frame2[19][1] = 3'h0;
    // frame2[19][2] = 3'h0;
    // frame2[19][3] = 3'h0;
    // frame2[19][4] = 3'h0;
    // frame2[19][5] = 3'h0;
    // frame2[19][6] = 3'h0;
    // frame2[19][7] = 3'h1;
    // frame2[19][8] = 3'h2;
    // frame2[19][9] = 3'h2;
    // frame2[19][10] = 3'h5;
    // frame2[19][11] = 3'h5;
    // frame2[19][12] = 3'h5;
    // frame2[19][13] = 3'h5;
    // frame2[19][14] = 3'h5;
    // frame2[19][15] = 3'h5;
    // frame2[19][16] = 3'h5;
    // frame2[19][17] = 3'h5;
    // frame2[19][18] = 3'h5;
    // frame2[19][19] = 3'h5;
    // frame2[19][20] = 3'h5;
    // frame2[19][21] = 3'h5;
    // frame2[19][22] = 3'h2;
    // frame2[19][23] = 3'h2;
    // frame2[19][24] = 3'h1;
    // frame2[19][25] = 3'h0;
    // frame2[19][26] = 3'h0;
    // frame2[19][27] = 3'h0;
    // frame2[19][28] = 3'h0;
    // frame2[19][29] = 3'h0;
    // frame2[19][30] = 3'h0;
    // frame2[19][31] = 3'h0;
    // frame2[20][0] = 3'h0;
    // frame2[20][1] = 3'h0;
    // frame2[20][2] = 3'h0;
    // frame2[20][3] = 3'h0;
    // frame2[20][4] = 3'h0;
    // frame2[20][5] = 3'h0;
    // frame2[20][6] = 3'h0;
    // frame2[20][7] = 3'h1;
    // frame2[20][8] = 3'h1;
    // frame2[20][9] = 3'h2;
    // frame2[20][10] = 3'h2;
    // frame2[20][11] = 3'h2;
    // frame2[20][12] = 3'h5;
    // frame2[20][13] = 3'h5;
    // frame2[20][14] = 3'h5;
    // frame2[20][15] = 3'h5;
    // frame2[20][16] = 3'h5;
    // frame2[20][17] = 3'h5;
    // frame2[20][18] = 3'h5;
    // frame2[20][19] = 3'h5;
    // frame2[20][20] = 3'h2;
    // frame2[20][21] = 3'h2;
    // frame2[20][22] = 3'h2;
    // frame2[20][23] = 3'h1;
    // frame2[20][24] = 3'h1;
    // frame2[20][25] = 3'h0;
    // frame2[20][26] = 3'h0;
    // frame2[20][27] = 3'h0;
    // frame2[20][28] = 3'h0;
    // frame2[20][29] = 3'h0;
    // frame2[20][30] = 3'h0;
    // frame2[20][31] = 3'h0;
    // frame2[21][0] = 3'h0;
    // frame2[21][1] = 3'h0;
    // frame2[21][2] = 3'h0;
    // frame2[21][3] = 3'h0;
    // frame2[21][4] = 3'h0;
    // frame2[21][5] = 3'h0;
    // frame2[21][6] = 3'h0;
    // frame2[21][7] = 3'h1;
    // frame2[21][8] = 3'h1;
    // frame2[21][9] = 3'h1;
    // frame2[21][10] = 3'h1;
    // frame2[21][11] = 3'h1;
    // frame2[21][12] = 3'h2;
    // frame2[21][13] = 3'h5;
    // frame2[21][14] = 3'h5;
    // frame2[21][15] = 3'h5;
    // frame2[21][16] = 3'h5;
    // frame2[21][17] = 3'h5;
    // frame2[21][18] = 3'h5;
    // frame2[21][19] = 3'h2;
    // frame2[21][20] = 3'h1;
    // frame2[21][21] = 3'h1;
    // frame2[21][22] = 3'h1;
    // frame2[21][23] = 3'h1;
    // frame2[21][24] = 3'h1;
    // frame2[21][25] = 3'h0;
    // frame2[21][26] = 3'h0;
    // frame2[21][27] = 3'h0;
    // frame2[21][28] = 3'h0;
    // frame2[21][29] = 3'h0;
    // frame2[21][30] = 3'h0;
    // frame2[21][31] = 3'h0;
    // frame2[22][0] = 3'h0;
    // frame2[22][1] = 3'h0;
    // frame2[22][2] = 3'h0;
    // frame2[22][3] = 3'h0;
    // frame2[22][4] = 3'h0;
    // frame2[22][5] = 3'h0;
    // frame2[22][6] = 3'h0;
    // frame2[22][7] = 3'h0;
    // frame2[22][8] = 3'h1;
    // frame2[22][9] = 3'h3;
    // frame2[22][10] = 3'h4;
    // frame2[22][11] = 3'h1;
    // frame2[22][12] = 3'h1;
    // frame2[22][13] = 3'h2;
    // frame2[22][14] = 3'h2;
    // frame2[22][15] = 3'h5;
    // frame2[22][16] = 3'h5;
    // frame2[22][17] = 3'h2;
    // frame2[22][18] = 3'h2;
    // frame2[22][19] = 3'h1;
    // frame2[22][20] = 3'h1;
    // frame2[22][21] = 3'h4;
    // frame2[22][22] = 3'h3;
    // frame2[22][23] = 3'h1;
    // frame2[22][24] = 3'h0;
    // frame2[22][25] = 3'h0;
    // frame2[22][26] = 3'h0;
    // frame2[22][27] = 3'h0;
    // frame2[22][28] = 3'h0;
    // frame2[22][29] = 3'h0;
    // frame2[22][30] = 3'h0;
    // frame2[22][31] = 3'h0;
    // frame2[23][0] = 3'h0;
    // frame2[23][1] = 3'h0;
    // frame2[23][2] = 3'h0;
    // frame2[23][3] = 3'h0;
    // frame2[23][4] = 3'h0;
    // frame2[23][5] = 3'h0;
    // frame2[23][6] = 3'h0;
    // frame2[23][7] = 3'h0;
    // frame2[23][8] = 3'h0;
    // frame2[23][9] = 3'h1;
    // frame2[23][10] = 3'h3;
    // frame2[23][11] = 3'h4;
    // frame2[23][12] = 3'h1;
    // frame2[23][13] = 3'h1;
    // frame2[23][14] = 3'h1;
    // frame2[23][15] = 3'h2;
    // frame2[23][16] = 3'h2;
    // frame2[23][17] = 3'h1;
    // frame2[23][18] = 3'h1;
    // frame2[23][19] = 3'h1;
    // frame2[23][20] = 3'h4;
    // frame2[23][21] = 3'h3;
    // frame2[23][22] = 3'h1;
    // frame2[23][23] = 3'h0;
    // frame2[23][24] = 3'h0;
    // frame2[23][25] = 3'h0;
    // frame2[23][26] = 3'h0;
    // frame2[23][27] = 3'h0;
    // frame2[23][28] = 3'h0;
    // frame2[23][29] = 3'h0;
    // frame2[23][30] = 3'h0;
    // frame2[23][31] = 3'h0;
    // frame2[24][0] = 3'h0;
    // frame2[24][1] = 3'h0;
    // frame2[24][2] = 3'h0;
    // frame2[24][3] = 3'h0;
    // frame2[24][4] = 3'h0;
    // frame2[24][5] = 3'h0;
    // frame2[24][6] = 3'h0;
    // frame2[24][7] = 3'h0;
    // frame2[24][8] = 3'h0;
    // frame2[24][9] = 3'h0;
    // frame2[24][10] = 3'h1;
    // frame2[24][11] = 3'h3;
    // frame2[24][12] = 3'h4;
    // frame2[24][13] = 3'h4;
    // frame2[24][14] = 3'h1;
    // frame2[24][15] = 3'h1;
    // frame2[24][16] = 3'h1;
    // frame2[24][17] = 3'h1;
    // frame2[24][18] = 3'h4;
    // frame2[24][19] = 3'h4;
    // frame2[24][20] = 3'h3;
    // frame2[24][21] = 3'h1;
    // frame2[24][22] = 3'h0;
    // frame2[24][23] = 3'h0;
    // frame2[24][24] = 3'h0;
    // frame2[24][25] = 3'h0;
    // frame2[24][26] = 3'h0;
    // frame2[24][27] = 3'h0;
    // frame2[24][28] = 3'h0;
    // frame2[24][29] = 3'h0;
    // frame2[24][30] = 3'h0;
    // frame2[24][31] = 3'h0;
    // frame2[25][0] = 3'h0;
    // frame2[25][1] = 3'h0;
    // frame2[25][2] = 3'h0;
    // frame2[25][3] = 3'h0;
    // frame2[25][4] = 3'h0;
    // frame2[25][5] = 3'h0;
    // frame2[25][6] = 3'h0;
    // frame2[25][7] = 3'h0;
    // frame2[25][8] = 3'h0;
    // frame2[25][9] = 3'h0;
    // frame2[25][10] = 3'h0;
    // frame2[25][11] = 3'h1;
    // frame2[25][12] = 3'h1;
    // frame2[25][13] = 3'h3;
    // frame2[25][14] = 3'h4;
    // frame2[25][15] = 3'h1;
    // frame2[25][16] = 3'h1;
    // frame2[25][17] = 3'h4;
    // frame2[25][18] = 3'h3;
    // frame2[25][19] = 3'h1;
    // frame2[25][20] = 3'h1;
    // frame2[25][21] = 3'h0;
    // frame2[25][22] = 3'h0;
    // frame2[25][23] = 3'h0;
    // frame2[25][24] = 3'h0;
    // frame2[25][25] = 3'h0;
    // frame2[25][26] = 3'h0;
    // frame2[25][27] = 3'h0;
    // frame2[25][28] = 3'h0;
    // frame2[25][29] = 3'h0;
    // frame2[25][30] = 3'h0;
    // frame2[25][31] = 3'h0;
    // frame2[26][0] = 3'h0;
    // frame2[26][1] = 3'h0;
    // frame2[26][2] = 3'h0;
    // frame2[26][3] = 3'h0;
    // frame2[26][4] = 3'h0;
    // frame2[26][5] = 3'h0;
    // frame2[26][6] = 3'h0;
    // frame2[26][7] = 3'h0;
    // frame2[26][8] = 3'h0;
    // frame2[26][9] = 3'h0;
    // frame2[26][10] = 3'h0;
    // frame2[26][11] = 3'h0;
    // frame2[26][12] = 3'h1;
    // frame2[26][13] = 3'h1;
    // frame2[26][14] = 3'h3;
    // frame2[26][15] = 3'h4;
    // frame2[26][16] = 3'h4;
    // frame2[26][17] = 3'h3;
    // frame2[26][18] = 3'h1;
    // frame2[26][19] = 3'h1;
    // frame2[26][20] = 3'h0;
    // frame2[26][21] = 3'h0;
    // frame2[26][22] = 3'h0;
    // frame2[26][23] = 3'h0;
    // frame2[26][24] = 3'h0;
    // frame2[26][25] = 3'h0;
    // frame2[26][26] = 3'h0;
    // frame2[26][27] = 3'h0;
    // frame2[26][28] = 3'h0;
    // frame2[26][29] = 3'h0;
    // frame2[26][30] = 3'h0;
    // frame2[26][31] = 3'h0;
    // frame2[27][0] = 3'h0;
    // frame2[27][1] = 3'h0;
    // frame2[27][2] = 3'h0;
    // frame2[27][3] = 3'h0;
    // frame2[27][4] = 3'h0;
    // frame2[27][5] = 3'h0;
    // frame2[27][6] = 3'h0;
    // frame2[27][7] = 3'h0;
    // frame2[27][8] = 3'h0;
    // frame2[27][9] = 3'h0;
    // frame2[27][10] = 3'h0;
    // frame2[27][11] = 3'h0;
    // frame2[27][12] = 3'h1;
    // frame2[27][13] = 3'h0;
    // frame2[27][14] = 3'h1;
    // frame2[27][15] = 3'h1;
    // frame2[27][16] = 3'h1;
    // frame2[27][17] = 3'h1;
    // frame2[27][18] = 3'h0;
    // frame2[27][19] = 3'h1;
    // frame2[27][20] = 3'h0;
    // frame2[27][21] = 3'h0;
    // frame2[27][22] = 3'h0;
    // frame2[27][23] = 3'h0;
    // frame2[27][24] = 3'h0;
    // frame2[27][25] = 3'h0;
    // frame2[27][26] = 3'h0;
    // frame2[27][27] = 3'h0;
    // frame2[27][28] = 3'h0;
    // frame2[27][29] = 3'h0;
    // frame2[27][30] = 3'h0;
    // frame2[27][31] = 3'h0;
    // frame2[28][0] = 3'h0;
    // frame2[28][1] = 3'h0;
    // frame2[28][2] = 3'h0;
    // frame2[28][3] = 3'h0;
    // frame2[28][4] = 3'h0;
    // frame2[28][5] = 3'h0;
    // frame2[28][6] = 3'h0;
    // frame2[28][7] = 3'h0;
    // frame2[28][8] = 3'h0;
    // frame2[28][9] = 3'h0;
    // frame2[28][10] = 3'h0;
    // frame2[28][11] = 3'h0;
    // frame2[28][12] = 3'h1;
    // frame2[28][13] = 3'h0;
    // frame2[28][14] = 3'h0;
    // frame2[28][15] = 3'h0;
    // frame2[28][16] = 3'h0;
    // frame2[28][17] = 3'h0;
    // frame2[28][18] = 3'h0;
    // frame2[28][19] = 3'h1;
    // frame2[28][20] = 3'h0;
    // frame2[28][21] = 3'h0;
    // frame2[28][22] = 3'h0;
    // frame2[28][23] = 3'h0;
    // frame2[28][24] = 3'h0;
    // frame2[28][25] = 3'h0;
    // frame2[28][26] = 3'h0;
    // frame2[28][27] = 3'h0;
    // frame2[28][28] = 3'h0;
    // frame2[28][29] = 3'h0;
    // frame2[28][30] = 3'h0;
    // frame2[28][31] = 3'h0;
    // frame2[29][0] = 3'h0;
    // frame2[29][1] = 3'h0;
    // frame2[29][2] = 3'h0;
    // frame2[29][3] = 3'h0;
    // frame2[29][4] = 3'h0;
    // frame2[29][5] = 3'h0;
    // frame2[29][6] = 3'h0;
    // frame2[29][7] = 3'h0;
    // frame2[29][8] = 3'h0;
    // frame2[29][9] = 3'h0;
    // frame2[29][10] = 3'h0;
    // frame2[29][11] = 3'h0;
    // frame2[29][12] = 3'h1;
    // frame2[29][13] = 3'h0;
    // frame2[29][14] = 3'h0;
    // frame2[29][15] = 3'h0;
    // frame2[29][16] = 3'h0;
    // frame2[29][17] = 3'h0;
    // frame2[29][18] = 3'h0;
    // frame2[29][19] = 3'h1;
    // frame2[29][20] = 3'h0;
    // frame2[29][21] = 3'h0;
    // frame2[29][22] = 3'h0;
    // frame2[29][23] = 3'h0;
    // frame2[29][24] = 3'h0;
    // frame2[29][25] = 3'h0;
    // frame2[29][26] = 3'h0;
    // frame2[29][27] = 3'h0;
    // frame2[29][28] = 3'h0;
    // frame2[29][29] = 3'h0;
    // frame2[29][30] = 3'h0;
    // frame2[29][31] = 3'h0;
    // frame2[30][0] = 3'h0;
    // frame2[30][1] = 3'h0;
    // frame2[30][2] = 3'h0;
    // frame2[30][3] = 3'h0;
    // frame2[30][4] = 3'h0;
    // frame2[30][5] = 3'h0;
    // frame2[30][6] = 3'h0;
    // frame2[30][7] = 3'h0;
    // frame2[30][8] = 3'h0;
    // frame2[30][9] = 3'h0;
    // frame2[30][10] = 3'h0;
    // frame2[30][11] = 3'h1;
    // frame2[30][12] = 3'h1;
    // frame2[30][13] = 3'h1;
    // frame2[30][14] = 3'h0;
    // frame2[30][15] = 3'h0;
    // frame2[30][16] = 3'h0;
    // frame2[30][17] = 3'h0;
    // frame2[30][18] = 3'h1;
    // frame2[30][19] = 3'h1;
    // frame2[30][20] = 3'h1;
    // frame2[30][21] = 3'h0;
    // frame2[30][22] = 3'h0;
    // frame2[30][23] = 3'h0;
    // frame2[30][24] = 3'h0;
    // frame2[30][25] = 3'h0;
    // frame2[30][26] = 3'h0;
    // frame2[30][27] = 3'h0;
    // frame2[30][28] = 3'h0;
    // frame2[30][29] = 3'h0;
    // frame2[30][30] = 3'h0;
    // frame2[30][31] = 3'h0;
    // frame2[31][0] = 3'h0;
    // frame2[31][1] = 3'h0;
    // frame2[31][2] = 3'h0;
    // frame2[31][3] = 3'h0;
    // frame2[31][4] = 3'h0;
    // frame2[31][5] = 3'h0;
    // frame2[31][6] = 3'h0;
    // frame2[31][7] = 3'h0;
    // frame2[31][8] = 3'h0;
    // frame2[31][9] = 3'h0;
    // frame2[31][10] = 3'h1;
    // frame2[31][11] = 3'h0;
    // frame2[31][12] = 3'h1;
    // frame2[31][13] = 3'h0;
    // frame2[31][14] = 3'h1;
    // frame2[31][15] = 3'h0;
    // frame2[31][16] = 3'h0;
    // frame2[31][17] = 3'h1;
    // frame2[31][18] = 3'h0;
    // frame2[31][19] = 3'h1;
    // frame2[31][20] = 3'h0;
    // frame2[31][21] = 3'h1;
    // frame2[31][22] = 3'h0;
    // frame2[31][23] = 3'h0;
    // frame2[31][24] = 3'h0;
    // frame2[31][25] = 3'h0;
    // frame2[31][26] = 3'h0;
    // frame2[31][27] = 3'h0;
    // frame2[31][28] = 3'h0;
    // frame2[31][29] = 3'h0;
    // frame2[31][30] = 3'h0;
    // frame2[31][31] = 3'h0;
end