reg [2:0] frame1 [0:24][0:24];
initial begin
    frame1[0][0] = 3'd0;
    frame1[0][1] = 3'd0;
    frame1[0][2] = 3'd0;
    frame1[0][3] = 3'd0;
    frame1[0][4] = 3'd0;
    frame1[0][5] = 3'd0;
    frame1[0][6] = 3'd0;
    frame1[0][7] = 3'd0;
    frame1[0][8] = 3'd0;
    frame1[0][9] = 3'd0;
    frame1[0][10] = 3'd0;
    frame1[0][11] = 3'd0;
    frame1[0][12] = 3'd0;
    frame1[0][13] = 3'd0;
    frame1[0][14] = 3'd0;
    frame1[0][15] = 3'd0;
    frame1[0][16] = 3'd0;
    frame1[0][17] = 3'd0;
    frame1[0][18] = 3'd0;
    frame1[0][19] = 3'd0;
    frame1[0][20] = 3'd0;
    frame1[0][21] = 3'd0;
    frame1[0][22] = 3'd0;
    frame1[0][23] = 3'd0;
    frame1[0][24] = 3'd0;
    frame1[1][0] = 3'd0;
    frame1[1][1] = 3'd0;
    frame1[1][2] = 3'd0;
    frame1[1][3] = 3'd0;
    frame1[1][4] = 3'd0;
    frame1[1][5] = 3'd1;
    frame1[1][6] = 3'd1;
    frame1[1][7] = 3'd1;
    frame1[1][8] = 3'd1;
    frame1[1][9] = 3'd0;
    frame1[1][10] = 3'd0;
    frame1[1][11] = 3'd0;
    frame1[1][12] = 3'd0;
    frame1[1][13] = 3'd0;
    frame1[1][14] = 3'd0;
    frame1[1][15] = 3'd0;
    frame1[1][16] = 3'd0;
    frame1[1][17] = 3'd0;
    frame1[1][18] = 3'd0;
    frame1[1][19] = 3'd0;
    frame1[1][20] = 3'd0;
    frame1[1][21] = 3'd0;
    frame1[1][22] = 3'd0;
    frame1[1][23] = 3'd0;
    frame1[1][24] = 3'd0;
    frame1[2][0] = 3'd0;
    frame1[2][1] = 3'd0;
    frame1[2][2] = 3'd0;
    frame1[2][3] = 3'd1;
    frame1[2][4] = 3'd1;
    frame1[2][5] = 3'd2;
    frame1[2][6] = 3'd2;
    frame1[2][7] = 3'd2;
    frame1[2][8] = 3'd2;
    frame1[2][9] = 3'd1;
    frame1[2][10] = 3'd0;
    frame1[2][11] = 3'd0;
    frame1[2][12] = 3'd0;
    frame1[2][13] = 3'd0;
    frame1[2][14] = 3'd0;
    frame1[2][15] = 3'd0;
    frame1[2][16] = 3'd0;
    frame1[2][17] = 3'd0;
    frame1[2][18] = 3'd0;
    frame1[2][19] = 3'd0;
    frame1[2][20] = 3'd0;
    frame1[2][21] = 3'd0;
    frame1[2][22] = 3'd0;
    frame1[2][23] = 3'd0;
    frame1[2][24] = 3'd0;
    frame1[3][0] = 3'd0;
    frame1[3][1] = 3'd0;
    frame1[3][2] = 3'd0;
    frame1[3][3] = 3'd1;
    frame1[3][4] = 3'd2;
    frame1[3][5] = 3'd1;
    frame1[3][6] = 3'd1;
    frame1[3][7] = 3'd2;
    frame1[3][8] = 3'd2;
    frame1[3][9] = 3'd1;
    frame1[3][10] = 3'd0;
    frame1[3][11] = 3'd0;
    frame1[3][12] = 3'd0;
    frame1[3][13] = 3'd0;
    frame1[3][14] = 3'd0;
    frame1[3][15] = 3'd0;
    frame1[3][16] = 3'd0;
    frame1[3][17] = 3'd0;
    frame1[3][18] = 3'd0;
    frame1[3][19] = 3'd0;
    frame1[3][20] = 3'd0;
    frame1[3][21] = 3'd0;
    frame1[3][22] = 3'd0;
    frame1[3][23] = 3'd0;
    frame1[3][24] = 3'd0;
    frame1[4][0] = 3'd0;
    frame1[4][1] = 3'd0;
    frame1[4][2] = 3'd0;
    frame1[4][3] = 3'd1;
    frame1[4][4] = 3'd2;
    frame1[4][5] = 3'd1;
    frame1[4][6] = 3'd2;
    frame1[4][7] = 3'd2;
    frame1[4][8] = 3'd2;
    frame1[4][9] = 3'd1;
    frame1[4][10] = 3'd0;
    frame1[4][11] = 3'd0;
    frame1[4][12] = 3'd0;
    frame1[4][13] = 3'd0;
    frame1[4][14] = 3'd0;
    frame1[4][15] = 3'd0;
    frame1[4][16] = 3'd0;
    frame1[4][17] = 3'd0;
    frame1[4][18] = 3'd0;
    frame1[4][19] = 3'd0;
    frame1[4][20] = 3'd0;
    frame1[4][21] = 3'd0;
    frame1[4][22] = 3'd0;
    frame1[4][23] = 3'd0;
    frame1[4][24] = 3'd0;
    frame1[5][0] = 3'd0;
    frame1[5][1] = 3'd1;
    frame1[5][2] = 3'd1;
    frame1[5][3] = 3'd1;
    frame1[5][4] = 3'd1;
    frame1[5][5] = 3'd2;
    frame1[5][6] = 3'd2;
    frame1[5][7] = 3'd2;
    frame1[5][8] = 3'd3;
    frame1[5][9] = 3'd1;
    frame1[5][10] = 3'd0;
    frame1[5][11] = 3'd0;
    frame1[5][12] = 3'd0;
    frame1[5][13] = 3'd0;
    frame1[5][14] = 3'd0;
    frame1[5][15] = 3'd0;
    frame1[5][16] = 3'd0;
    frame1[5][17] = 3'd0;
    frame1[5][18] = 3'd0;
    frame1[5][19] = 3'd0;
    frame1[5][20] = 3'd0;
    frame1[5][21] = 3'd0;
    frame1[5][22] = 3'd0;
    frame1[5][23] = 3'd0;
    frame1[5][24] = 3'd0;
    frame1[6][0] = 3'd0;
    frame1[6][1] = 3'd0;
    frame1[6][2] = 3'd0;
    frame1[6][3] = 3'd0;
    frame1[6][4] = 3'd0;
    frame1[6][5] = 3'd1;
    frame1[6][6] = 3'd1;
    frame1[6][7] = 3'd3;
    frame1[6][8] = 3'd3;
    frame1[6][9] = 3'd1;
    frame1[6][10] = 3'd0;
    frame1[6][11] = 3'd0;
    frame1[6][12] = 3'd0;
    frame1[6][13] = 3'd0;
    frame1[6][14] = 3'd0;
    frame1[6][15] = 3'd0;
    frame1[6][16] = 3'd0;
    frame1[6][17] = 3'd0;
    frame1[6][18] = 3'd0;
    frame1[6][19] = 3'd0;
    frame1[6][20] = 3'd0;
    frame1[6][21] = 3'd0;
    frame1[6][22] = 3'd0;
    frame1[6][23] = 3'd0;
    frame1[6][24] = 3'd0;
    frame1[7][0] = 3'd0;
    frame1[7][1] = 3'd0;
    frame1[7][2] = 3'd0;
    frame1[7][3] = 3'd0;
    frame1[7][4] = 3'd0;
    frame1[7][5] = 3'd0;
    frame1[7][6] = 3'd1;
    frame1[7][7] = 3'd3;
    frame1[7][8] = 3'd2;
    frame1[7][9] = 3'd1;
    frame1[7][10] = 3'd0;
    frame1[7][11] = 3'd0;
    frame1[7][12] = 3'd0;
    frame1[7][13] = 3'd0;
    frame1[7][14] = 3'd0;
    frame1[7][15] = 3'd0;
    frame1[7][16] = 3'd0;
    frame1[7][17] = 3'd0;
    frame1[7][18] = 3'd0;
    frame1[7][19] = 3'd0;
    frame1[7][20] = 3'd0;
    frame1[7][21] = 3'd0;
    frame1[7][22] = 3'd0;
    frame1[7][23] = 3'd0;
    frame1[7][24] = 3'd0;
    frame1[8][0] = 3'd0;
    frame1[8][1] = 3'd0;
    frame1[8][2] = 3'd0;
    frame1[8][3] = 3'd0;
    frame1[8][4] = 3'd0;
    frame1[8][5] = 3'd0;
    frame1[8][6] = 3'd1;
    frame1[8][7] = 3'd2;
    frame1[8][8] = 3'd2;
    frame1[8][9] = 3'd1;
    frame1[8][10] = 3'd0;
    frame1[8][11] = 3'd0;
    frame1[8][12] = 3'd0;
    frame1[8][13] = 3'd0;
    frame1[8][14] = 3'd0;
    frame1[8][15] = 3'd0;
    frame1[8][16] = 3'd0;
    frame1[8][17] = 3'd0;
    frame1[8][18] = 3'd0;
    frame1[8][19] = 3'd0;
    frame1[8][20] = 3'd0;
    frame1[8][21] = 3'd0;
    frame1[8][22] = 3'd0;
    frame1[8][23] = 3'd0;
    frame1[8][24] = 3'd0;
    frame1[9][0] = 3'd0;
    frame1[9][1] = 3'd0;
    frame1[9][2] = 3'd0;
    frame1[9][3] = 3'd0;
    frame1[9][4] = 3'd0;
    frame1[9][5] = 3'd0;
    frame1[9][6] = 3'd1;
    frame1[9][7] = 3'd2;
    frame1[9][8] = 3'd2;
    frame1[9][9] = 3'd1;
    frame1[9][10] = 3'd0;
    frame1[9][11] = 3'd0;
    frame1[9][12] = 3'd0;
    frame1[9][13] = 3'd0;
    frame1[9][14] = 3'd0;
    frame1[9][15] = 3'd0;
    frame1[9][16] = 3'd0;
    frame1[9][17] = 3'd0;
    frame1[9][18] = 3'd0;
    frame1[9][19] = 3'd0;
    frame1[9][20] = 3'd0;
    frame1[9][21] = 3'd0;
    frame1[9][22] = 3'd0;
    frame1[9][23] = 3'd0;
    frame1[9][24] = 3'd0;
    frame1[10][0] = 3'd0;
    frame1[10][1] = 3'd0;
    frame1[10][2] = 3'd0;
    frame1[10][3] = 3'd0;
    frame1[10][4] = 3'd0;
    frame1[10][5] = 3'd0;
    frame1[10][6] = 3'd1;
    frame1[10][7] = 3'd2;
    frame1[10][8] = 3'd2;
    frame1[10][9] = 3'd1;
    frame1[10][10] = 3'd0;
    frame1[10][11] = 3'd0;
    frame1[10][12] = 3'd0;
    frame1[10][13] = 3'd0;
    frame1[10][14] = 3'd0;
    frame1[10][15] = 3'd0;
    frame1[10][16] = 3'd0;
    frame1[10][17] = 3'd0;
    frame1[10][18] = 3'd0;
    frame1[10][19] = 3'd0;
    frame1[10][20] = 3'd0;
    frame1[10][21] = 3'd0;
    frame1[10][22] = 3'd0;
    frame1[10][23] = 3'd0;
    frame1[10][24] = 3'd0;
    frame1[11][0] = 3'd0;
    frame1[11][1] = 3'd0;
    frame1[11][2] = 3'd0;
    frame1[11][3] = 3'd0;
    frame1[11][4] = 3'd0;
    frame1[11][5] = 3'd1;
    frame1[11][6] = 3'd1;
    frame1[11][7] = 3'd2;
    frame1[11][8] = 3'd2;
    frame1[11][9] = 3'd1;
    frame1[11][10] = 3'd1;
    frame1[11][11] = 3'd0;
    frame1[11][12] = 3'd0;
    frame1[11][13] = 3'd0;
    frame1[11][14] = 3'd0;
    frame1[11][15] = 3'd0;
    frame1[11][16] = 3'd0;
    frame1[11][17] = 3'd0;
    frame1[11][18] = 3'd0;
    frame1[11][19] = 3'd0;
    frame1[11][20] = 3'd0;
    frame1[11][21] = 3'd0;
    frame1[11][22] = 3'd0;
    frame1[11][23] = 3'd0;
    frame1[11][24] = 3'd0;
    frame1[12][0] = 3'd0;
    frame1[12][1] = 3'd0;
    frame1[12][2] = 3'd0;
    frame1[12][3] = 3'd0;
    frame1[12][4] = 3'd0;
    frame1[12][5] = 3'd1;
    frame1[12][6] = 3'd4;
    frame1[12][7] = 3'd4;
    frame1[12][8] = 3'd4;
    frame1[12][9] = 3'd2;
    frame1[12][10] = 3'd1;
    frame1[12][11] = 3'd1;
    frame1[12][12] = 3'd1;
    frame1[12][13] = 3'd1;
    frame1[12][14] = 3'd1;
    frame1[12][15] = 3'd1;
    frame1[12][16] = 3'd0;
    frame1[12][17] = 3'd0;
    frame1[12][18] = 3'd0;
    frame1[12][19] = 3'd0;
    frame1[12][20] = 3'd0;
    frame1[12][21] = 3'd0;
    frame1[12][22] = 3'd1;
    frame1[12][23] = 3'd1;
    frame1[12][24] = 3'd0;
    frame1[13][0] = 3'd0;
    frame1[13][1] = 3'd0;
    frame1[13][2] = 3'd0;
    frame1[13][3] = 3'd1;
    frame1[13][4] = 3'd1;
    frame1[13][5] = 3'd4;
    frame1[13][6] = 3'd4;
    frame1[13][7] = 3'd5;
    frame1[13][8] = 3'd5;
    frame1[13][9] = 3'd5;
    frame1[13][10] = 3'd5;
    frame1[13][11] = 3'd5;
    frame1[13][12] = 3'd5;
    frame1[13][13] = 3'd5;
    frame1[13][14] = 3'd5;
    frame1[13][15] = 3'd5;
    frame1[13][16] = 3'd5;
    frame1[13][17] = 3'd5;
    frame1[13][18] = 3'd1;
    frame1[13][19] = 3'd1;
    frame1[13][20] = 3'd1;
    frame1[13][21] = 3'd5;
    frame1[13][22] = 3'd5;
    frame1[13][23] = 3'd1;
    frame1[13][24] = 3'd0;
    frame1[14][0] = 3'd0;
    frame1[14][1] = 3'd0;
    frame1[14][2] = 3'd0;
    frame1[14][3] = 3'd1;
    frame1[14][4] = 3'd4;
    frame1[14][5] = 3'd4;
    frame1[14][6] = 3'd5;
    frame1[14][7] = 3'd5;
    frame1[14][8] = 3'd5;
    frame1[14][9] = 3'd5;
    frame1[14][10] = 3'd2;
    frame1[14][11] = 3'd2;
    frame1[14][12] = 3'd5;
    frame1[14][13] = 3'd5;
    frame1[14][14] = 3'd5;
    frame1[14][15] = 3'd5;
    frame1[14][16] = 3'd5;
    frame1[14][17] = 3'd5;
    frame1[14][18] = 3'd5;
    frame1[14][19] = 3'd5;
    frame1[14][20] = 3'd5;
    frame1[14][21] = 3'd5;
    frame1[14][22] = 3'd5;
    frame1[14][23] = 3'd1;
    frame1[14][24] = 3'd0;
    frame1[15][0] = 3'd0;
    frame1[15][1] = 3'd0;
    frame1[15][2] = 3'd0;
    frame1[15][3] = 3'd1;
    frame1[15][4] = 3'd4;
    frame1[15][5] = 3'd4;
    frame1[15][6] = 3'd5;
    frame1[15][7] = 3'd5;
    frame1[15][8] = 3'd5;
    frame1[15][9] = 3'd5;
    frame1[15][10] = 3'd1;
    frame1[15][11] = 3'd2;
    frame1[15][12] = 3'd2;
    frame1[15][13] = 3'd5;
    frame1[15][14] = 3'd5;
    frame1[15][15] = 3'd5;
    frame1[15][16] = 3'd5;
    frame1[15][17] = 3'd5;
    frame1[15][18] = 3'd5;
    frame1[15][19] = 3'd5;
    frame1[15][20] = 3'd5;
    frame1[15][21] = 3'd5;
    frame1[15][22] = 3'd5;
    frame1[15][23] = 3'd1;
    frame1[15][24] = 3'd0;
    frame1[16][0] = 3'd0;
    frame1[16][1] = 3'd0;
    frame1[16][2] = 3'd0;
    frame1[16][3] = 3'd1;
    frame1[16][4] = 3'd4;
    frame1[16][5] = 3'd4;
    frame1[16][6] = 3'd4;
    frame1[16][7] = 3'd5;
    frame1[16][8] = 3'd5;
    frame1[16][9] = 3'd5;
    frame1[16][10] = 3'd5;
    frame1[16][11] = 3'd5;
    frame1[16][12] = 3'd5;
    frame1[16][13] = 3'd2;
    frame1[16][14] = 3'd2;
    frame1[16][15] = 3'd2;
    frame1[16][16] = 3'd2;
    frame1[16][17] = 3'd2;
    frame1[16][18] = 3'd2;
    frame1[16][19] = 3'd2;
    frame1[16][20] = 3'd3;
    frame1[16][21] = 3'd1;
    frame1[16][22] = 3'd1;
    frame1[16][23] = 3'd0;
    frame1[16][24] = 3'd0;
    frame1[17][0] = 3'd0;
    frame1[17][1] = 3'd0;
    frame1[17][2] = 3'd0;
    frame1[17][3] = 3'd1;
    frame1[17][4] = 3'd1;
    frame1[17][5] = 3'd4;
    frame1[17][6] = 3'd4;
    frame1[17][7] = 3'd4;
    frame1[17][8] = 3'd5;
    frame1[17][9] = 3'd5;
    frame1[17][10] = 3'd5;
    frame1[17][11] = 3'd5;
    frame1[17][12] = 3'd5;
    frame1[17][13] = 3'd1;
    frame1[17][14] = 3'd1;
    frame1[17][15] = 3'd1;
    frame1[17][16] = 3'd1;
    frame1[17][17] = 3'd1;
    frame1[17][18] = 3'd1;
    frame1[17][19] = 3'd1;
    frame1[17][20] = 3'd1;
    frame1[17][21] = 3'd1;
    frame1[17][22] = 3'd0;
    frame1[17][23] = 3'd0;
    frame1[17][24] = 3'd0;
    frame1[18][0] = 3'd0;
    frame1[18][1] = 3'd0;
    frame1[18][2] = 3'd0;
    frame1[18][3] = 3'd0;
    frame1[18][4] = 3'd0;
    frame1[18][5] = 3'd1;
    frame1[18][6] = 3'd4;
    frame1[18][7] = 3'd4;
    frame1[18][8] = 3'd4;
    frame1[18][9] = 3'd5;
    frame1[18][10] = 3'd5;
    frame1[18][11] = 3'd5;
    frame1[18][12] = 3'd5;
    frame1[18][13] = 3'd3;
    frame1[18][14] = 3'd3;
    frame1[18][15] = 3'd3;
    frame1[18][16] = 3'd3;
    frame1[18][17] = 3'd3;
    frame1[18][18] = 3'd3;
    frame1[18][19] = 3'd3;
    frame1[18][20] = 3'd1;
    frame1[18][21] = 3'd0;
    frame1[18][22] = 3'd0;
    frame1[18][23] = 3'd0;
    frame1[18][24] = 3'd0;
    frame1[19][0] = 3'd0;
    frame1[19][1] = 3'd0;
    frame1[19][2] = 3'd0;
    frame1[19][3] = 3'd0;
    frame1[19][4] = 3'd0;
    frame1[19][5] = 3'd1;
    frame1[19][6] = 3'd1;
    frame1[19][7] = 3'd4;
    frame1[19][8] = 3'd4;
    frame1[19][9] = 3'd4;
    frame1[19][10] = 3'd4;
    frame1[19][11] = 3'd4;
    frame1[19][12] = 3'd4;
    frame1[19][13] = 3'd4;
    frame1[19][14] = 3'd3;
    frame1[19][15] = 3'd3;
    frame1[19][16] = 3'd3;
    frame1[19][17] = 3'd4;
    frame1[19][18] = 3'd4;
    frame1[19][19] = 3'd1;
    frame1[19][20] = 3'd0;
    frame1[19][21] = 3'd0;
    frame1[19][22] = 3'd0;
    frame1[19][23] = 3'd0;
    frame1[19][24] = 3'd0;
    frame1[20][0] = 3'd0;
    frame1[20][1] = 3'd0;
    frame1[20][2] = 3'd0;
    frame1[20][3] = 3'd0;
    frame1[20][4] = 3'd0;
    frame1[20][5] = 3'd0;
    frame1[20][6] = 3'd0;
    frame1[20][7] = 3'd0;
    frame1[20][8] = 3'd1;
    frame1[20][9] = 3'd1;
    frame1[20][10] = 3'd1;
    frame1[20][11] = 3'd5;
    frame1[20][12] = 3'd5;
    frame1[20][13] = 3'd1;
    frame1[20][14] = 3'd1;
    frame1[20][15] = 3'd1;
    frame1[20][16] = 3'd1;
    frame1[20][17] = 3'd1;
    frame1[20][18] = 3'd0;
    frame1[20][19] = 3'd0;
    frame1[20][20] = 3'd0;
    frame1[20][21] = 3'd0;
    frame1[20][22] = 3'd0;
    frame1[20][23] = 3'd0;
    frame1[20][24] = 3'd0;
    frame1[21][0] = 3'd0;
    frame1[21][1] = 3'd0;
    frame1[21][2] = 3'd0;
    frame1[21][3] = 3'd0;
    frame1[21][4] = 3'd0;
    frame1[21][5] = 3'd0;
    frame1[21][6] = 3'd0;
    frame1[21][7] = 3'd0;
    frame1[21][8] = 3'd0;
    frame1[21][9] = 3'd0;
    frame1[21][10] = 3'd1;
    frame1[21][11] = 3'd1;
    frame1[21][12] = 3'd1;
    frame1[21][13] = 3'd1;
    frame1[21][14] = 3'd0;
    frame1[21][15] = 3'd1;
    frame1[21][16] = 3'd0;
    frame1[21][17] = 3'd0;
    frame1[21][18] = 3'd0;
    frame1[21][19] = 3'd0;
    frame1[21][20] = 3'd0;
    frame1[21][21] = 3'd0;
    frame1[21][22] = 3'd0;
    frame1[21][23] = 3'd0;
    frame1[21][24] = 3'd0;
    frame1[22][0] = 3'd0;
    frame1[22][1] = 3'd0;
    frame1[22][2] = 3'd0;
    frame1[22][3] = 3'd0;
    frame1[22][4] = 3'd0;
    frame1[22][5] = 3'd0;
    frame1[22][6] = 3'd0;
    frame1[22][7] = 3'd0;
    frame1[22][8] = 3'd0;
    frame1[22][9] = 3'd0;
    frame1[22][10] = 3'd0;
    frame1[22][11] = 3'd0;
    frame1[22][12] = 3'd1;
    frame1[22][13] = 3'd0;
    frame1[22][14] = 3'd0;
    frame1[22][15] = 3'd1;
    frame1[22][16] = 3'd0;
    frame1[22][17] = 3'd0;
    frame1[22][18] = 3'd0;
    frame1[22][19] = 3'd0;
    frame1[22][20] = 3'd0;
    frame1[22][21] = 3'd0;
    frame1[22][22] = 3'd0;
    frame1[22][23] = 3'd0;
    frame1[22][24] = 3'd0;
    frame1[23][0] = 3'd0;
    frame1[23][1] = 3'd0;
    frame1[23][2] = 3'd0;
    frame1[23][3] = 3'd0;
    frame1[23][4] = 3'd0;
    frame1[23][5] = 3'd0;
    frame1[23][6] = 3'd0;
    frame1[23][7] = 3'd0;
    frame1[23][8] = 3'd0;
    frame1[23][9] = 3'd0;
    frame1[23][10] = 3'd1;
    frame1[23][11] = 3'd1;
    frame1[23][12] = 3'd1;
    frame1[23][13] = 3'd0;
    frame1[23][14] = 3'd1;
    frame1[23][15] = 3'd1;
    frame1[23][16] = 3'd0;
    frame1[23][17] = 3'd0;
    frame1[23][18] = 3'd0;
    frame1[23][19] = 3'd0;
    frame1[23][20] = 3'd0;
    frame1[23][21] = 3'd0;
    frame1[23][22] = 3'd0;
    frame1[23][23] = 3'd0;
    frame1[23][24] = 3'd0;
    frame1[24][0] = 3'd0;
    frame1[24][1] = 3'd0;
    frame1[24][2] = 3'd0;
    frame1[24][3] = 3'd0;
    frame1[24][4] = 3'd0;
    frame1[24][5] = 3'd0;
    frame1[24][6] = 3'd0;
    frame1[24][7] = 3'd0;
    frame1[24][8] = 3'd0;
    frame1[24][9] = 3'd1;
    frame1[24][10] = 3'd1;
    frame1[24][11] = 3'd1;
    frame1[24][12] = 3'd1;
    frame1[24][13] = 3'd1;
    frame1[24][14] = 3'd1;
    frame1[24][15] = 3'd1;
    frame1[24][16] = 3'd0;
    frame1[24][17] = 3'd0;
    frame1[24][18] = 3'd0;
    frame1[24][19] = 3'd0;
    frame1[24][20] = 3'd0;
    frame1[24][21] = 3'd0;
    frame1[24][22] = 3'd0;
    frame1[24][23] = 3'd0;
    frame1[24][24] = 3'd0;
end