reg [5:0] frame3[7:0][31:0];
initial begin
    frame3[0][0] = 6'd0;
    frame3[1][0] = 6'd0;
    frame3[2][0] = 6'd0;
    frame3[3][0] = 6'd0;
    frame3[4][0] = 6'd0;
    frame3[5][0] = 6'd0;
    frame3[6][0] = 6'd0;
    frame3[7][0] = 6'd0;
    frame3[0][1] = 6'd0;
    frame3[1][1] = 6'd0;
    frame3[2][1] = 6'd0;
    frame3[3][1] = 6'd0;
    frame3[4][1] = 6'd0;
    frame3[5][1] = 6'd0;
    frame3[6][1] = 6'd0;
    frame3[7][1] = 6'd0;
    frame3[0][2] = 6'd0;
    frame3[1][2] = 6'd0;
    frame3[2][2] = 6'd0;
    frame3[3][2] = 6'd0;
    frame3[4][2] = 6'd0;
    frame3[5][2] = 6'd5;
    frame3[6][2] = 6'd2;
    frame3[7][2] = 6'd0;
    frame3[0][3] = 6'd0;
    frame3[1][3] = 6'd0;
    frame3[2][3] = 6'd0;
    frame3[3][3] = 6'd0;
    frame3[4][3] = 6'd0;
    frame3[5][3] = 6'd1;
    frame3[6][3] = 6'd8;
    frame3[7][3] = 6'd0;
    frame3[0][4] = 6'd0;
    frame3[1][4] = 6'd0;
    frame3[2][4] = 6'd0;
    frame3[3][4] = 6'd0;
    frame3[4][4] = 6'd0;
    frame3[5][4] = 6'd4;
    frame3[6][4] = 6'd13;
    frame3[7][4] = 6'd0;
    frame3[0][5] = 6'd0;
    frame3[1][5] = 6'd0;
    frame3[2][5] = 6'd0;
    frame3[3][5] = 6'd0;
    frame3[4][5] = 6'd0;
    frame3[5][5] = 6'd1;
    frame3[6][5] = 6'd13;
    frame3[7][5] = 6'd0;
    frame3[0][6] = 6'd0;
    frame3[1][6] = 6'd0;
    frame3[2][6] = 6'd0;
    frame3[3][6] = 6'd0;
    frame3[4][6] = 6'd0;
    frame3[5][6] = 6'd54;
    frame3[6][6] = 6'd4;
    frame3[7][6] = 6'd0;
    frame3[0][7] = 6'd0;
    frame3[1][7] = 6'd0;
    frame3[2][7] = 6'd0;
    frame3[3][7] = 6'd0;
    frame3[4][7] = 6'd0;
    frame3[5][7] = 6'd57;
    frame3[6][7] = 6'd8;
    frame3[7][7] = 6'd0;
    frame3[0][8] = 6'd0;
    frame3[1][8] = 6'd0;
    frame3[2][8] = 6'd0;
    frame3[3][8] = 6'd0;
    frame3[4][8] = 6'd0;
    frame3[5][8] = 6'd41;
    frame3[6][8] = 6'd0;
    frame3[7][8] = 6'd0;
    frame3[0][9] = 6'd0;
    frame3[1][9] = 6'd0;
    frame3[2][9] = 6'd0;
    frame3[3][9] = 6'd0;
    frame3[4][9] = 6'd0;
    frame3[5][9] = 6'd33;
    frame3[6][9] = 6'd0;
    frame3[7][9] = 6'd0;
    frame3[0][10] = 6'd0;
    frame3[1][10] = 6'd0;
    frame3[2][10] = 6'd0;
    frame3[3][10] = 6'd0;
    frame3[4][10] = 6'd0;
    frame3[5][10] = 6'd4;
    frame3[6][10] = 6'd0;
    frame3[7][10] = 6'd0;
    frame3[0][11] = 6'd0;
    frame3[1][11] = 6'd0;
    frame3[2][11] = 6'd0;
    frame3[3][11] = 6'd0;
    frame3[4][11] = 6'd0;
    frame3[5][11] = 6'd4;
    frame3[6][11] = 6'd0;
    frame3[7][11] = 6'd0;
    frame3[0][12] = 6'd0;
    frame3[1][12] = 6'd0;
    frame3[2][12] = 6'd0;
    frame3[3][12] = 6'd0;
    frame3[4][12] = 6'd0;
    frame3[5][12] = 6'd4;
    frame3[6][12] = 6'd0;
    frame3[7][12] = 6'd0;
    frame3[0][13] = 6'd0;
    frame3[1][13] = 6'd0;
    frame3[2][13] = 6'd0;
    frame3[3][13] = 6'd0;
    frame3[4][13] = 6'd0;
    frame3[5][13] = 6'd4;
    frame3[6][13] = 6'd0;
    frame3[7][13] = 6'd0;
    frame3[0][14] = 6'd0;
    frame3[1][14] = 6'd0;
    frame3[2][14] = 6'd0;
    frame3[3][14] = 6'd0;
    frame3[4][14] = 6'd0;
    frame3[5][14] = 6'd4;
    frame3[6][14] = 6'd0;
    frame3[7][14] = 6'd0;
    frame3[0][15] = 6'd0;
    frame3[1][15] = 6'd0;
    frame3[2][15] = 6'd0;
    frame3[3][15] = 6'd0;
    frame3[4][15] = 6'd3;
    frame3[5][15] = 6'd17;
    frame3[6][15] = 6'd0;
    frame3[7][15] = 6'd0;
    frame3[0][16] = 6'd49;
    frame3[1][16] = 6'd0;
    frame3[2][16] = 6'd0;
    frame3[3][16] = 6'd5;
    frame3[4][16] = 6'd1;
    frame3[5][16] = 6'd14;
    frame3[6][16] = 6'd11;
    frame3[7][16] = 6'd0;
    frame3[0][17] = 6'd7;
    frame3[1][17] = 6'd2;
    frame3[2][17] = 6'd5;
    frame3[3][17] = 6'd1;
    frame3[4][17] = 6'd1;
    frame3[5][17] = 6'd34;
    frame3[6][17] = 6'd29;
    frame3[7][17] = 6'd0;
    frame3[0][18] = 6'd7;
    frame3[1][18] = 6'd1;
    frame3[2][18] = 6'd1;
    frame3[3][18] = 6'd1;
    frame3[4][18] = 6'd1;
    frame3[5][18] = 6'd1;
    frame3[6][18] = 6'd10;
    frame3[7][18] = 6'd0;
    frame3[0][19] = 6'd3;
    frame3[1][19] = 6'd1;
    frame3[2][19] = 6'd1;
    frame3[3][19] = 6'd1;
    frame3[4][19] = 6'd18;
    frame3[5][19] = 6'd1;
    frame3[6][19] = 6'd10;
    frame3[7][19] = 6'd0;
    frame3[0][20] = 6'd0;
    frame3[1][20] = 6'd19;
    frame3[2][20] = 6'd1;
    frame3[3][20] = 6'd1;
    frame3[4][20] = 6'd7;
    frame3[5][20] = 6'd1;
    frame3[6][20] = 6'd10;
    frame3[7][20] = 6'd0;
    frame3[0][21] = 6'd0;
    frame3[1][21] = 6'd40;
    frame3[2][21] = 6'd1;
    frame3[3][21] = 6'd4;
    frame3[4][21] = 6'd1;
    frame3[5][21] = 6'd34;
    frame3[6][21] = 6'd10;
    frame3[7][21] = 6'd0;
    frame3[0][22] = 6'd0;
    frame3[1][22] = 6'd32;
    frame3[2][22] = 6'd0;
    frame3[3][22] = 6'd3;
    frame3[4][22] = 6'd1;
    frame3[5][22] = 6'd14;
    frame3[6][22] = 6'd11;
    frame3[7][22] = 6'd0;
    frame3[0][23] = 6'd0;
    frame3[1][23] = 6'd50;
    frame3[2][23] = 6'd20;
    frame3[3][23] = 6'd59;
    frame3[4][23] = 6'd1;
    frame3[5][23] = 6'd17;
    frame3[6][23] = 6'd0;
    frame3[7][23] = 6'd0;
    frame3[0][24] = 6'd0;
    frame3[1][24] = 6'd0;
    frame3[2][24] = 6'd25;
    frame3[3][24] = 6'd21;
    frame3[4][24] = 6'd6;
    frame3[5][24] = 6'd10;
    frame3[6][24] = 6'd0;
    frame3[7][24] = 6'd0;
    frame3[0][25] = 6'd0;
    frame3[1][25] = 6'd0;
    frame3[2][25] = 6'd26;
    frame3[3][25] = 6'd6;
    frame3[4][25] = 6'd6;
    frame3[5][25] = 6'd11;
    frame3[6][25] = 6'd0;
    frame3[7][25] = 6'd0;
    frame3[0][26] = 6'd0;
    frame3[1][26] = 6'd0;
    frame3[2][26] = 6'd0;
    frame3[3][26] = 6'd3;
    frame3[4][26] = 6'd8;
    frame3[5][26] = 6'd0;
    frame3[6][26] = 6'd0;
    frame3[7][26] = 6'd0;
    frame3[0][27] = 6'd0;
    frame3[1][27] = 6'd0;
    frame3[2][27] = 6'd0;
    frame3[3][27] = 6'd0;
    frame3[4][27] = 6'd0;
    frame3[5][27] = 6'd0;
    frame3[6][27] = 6'd0;
    frame3[7][27] = 6'd0;
    frame3[0][28] = 6'd0;
    frame3[1][28] = 6'd0;
    frame3[2][28] = 6'd0;
    frame3[3][28] = 6'd0;
    frame3[4][28] = 6'd0;
    frame3[5][28] = 6'd0;
    frame3[6][28] = 6'd0;
    frame3[7][28] = 6'd0;
    frame3[0][29] = 6'd0;
    frame3[1][29] = 6'd0;
    frame3[2][29] = 6'd0;
    frame3[3][29] = 6'd0;
    frame3[4][29] = 6'd0;
    frame3[5][29] = 6'd0;
    frame3[6][29] = 6'd0;
    frame3[7][29] = 6'd0;
    frame3[0][30] = 6'd0;
    frame3[1][30] = 6'd0;
    frame3[2][30] = 6'd0;
    frame3[3][30] = 6'd0;
    frame3[4][30] = 6'd0;
    frame3[5][30] = 6'd0;
    frame3[6][30] = 6'd0;
    frame3[7][30] = 6'd0;
    frame3[0][31] = 6'd0;
    frame3[1][31] = 6'd0;
    frame3[2][31] = 6'd0;
    frame3[3][31] = 6'd0;
    frame3[4][31] = 6'd0;
    frame3[5][31] = 6'd0;
    frame3[6][31] = 6'd0;
    frame3[7][31] = 6'd0;
end