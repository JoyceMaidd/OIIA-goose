reg [2:0] frame1 [0:15][0:15];
initial begin
    frame1[0][0] = 3'h0;
    frame1[0][1] = 3'h0;
    frame1[0][2] = 3'h0;
    frame1[0][3] = 3'h0;
    frame1[0][4] = 3'h0;
    frame1[0][5] = 3'h0;
    frame1[0][6] = 3'h0;
    frame1[0][7] = 3'h0;
    frame1[0][8] = 3'h0;
    frame1[0][9] = 3'h0;
    frame1[0][10] = 3'h0;
    frame1[0][11] = 3'h0;
    frame1[0][12] = 3'h0;
    frame1[0][13] = 3'h0;
    frame1[0][14] = 3'h0;
    frame1[0][15] = 3'h0;
    frame1[0][16] = 3'h0;
    frame1[0][17] = 3'h0;
    frame1[0][18] = 3'h0;
    frame1[0][19] = 3'h0;
    frame1[0][20] = 3'h0;
    frame1[0][21] = 3'h0;
    frame1[0][22] = 3'h0;
    frame1[0][23] = 3'h0;
    frame1[0][24] = 3'h0;
    // frame1[0][25] = 3'h0;
    // frame1[0][26] = 3'h0;
    // frame1[0][27] = 3'h0;
    // frame1[0][28] = 3'h0;
    // frame1[0][29] = 3'h0;
    // frame1[0][30] = 3'h0;
    // frame1[0][31] = 3'h0;
    frame1[1][0] = 3'h0;
    frame1[1][1] = 3'h0;
    frame1[1][2] = 3'h0;
    frame1[1][3] = 3'h0;
    frame1[1][4] = 3'h0;
    frame1[1][5] = 3'h0;
    frame1[1][6] = 3'h1;
    frame1[1][7] = 3'h1;
    frame1[1][8] = 3'h1;
    frame1[1][9] = 3'h1;
    frame1[1][10] = 3'h1;
    frame1[1][11] = 3'h1;
    frame1[1][12] = 3'h0;
    frame1[1][13] = 3'h0;
    frame1[1][14] = 3'h0;
    frame1[1][15] = 3'h0;
    frame1[1][16] = 3'h0;
    frame1[1][17] = 3'h0;
    frame1[1][18] = 3'h0;
    frame1[1][19] = 3'h0;
    frame1[1][20] = 3'h0;
    frame1[1][21] = 3'h0;
    frame1[1][22] = 3'h0;
    frame1[1][23] = 3'h0;
    frame1[1][24] = 3'h0;
    // frame1[1][25] = 3'h0;
    // frame1[1][26] = 3'h0;
    // frame1[1][27] = 3'h0;
    // frame1[1][28] = 3'h0;
    // frame1[1][29] = 3'h0;
    // frame1[1][30] = 3'h0;
    // frame1[1][31] = 3'h0;
    frame1[2][0] = 3'h0;
    frame1[2][1] = 3'h0;
    frame1[2][2] = 3'h0;
    frame1[2][3] = 3'h0;
    frame1[2][4] = 3'h0;
    frame1[2][5] = 3'h1;
    frame1[2][6] = 3'h1;
    frame1[2][7] = 3'h2;
    frame1[2][8] = 3'h2;
    frame1[2][9] = 3'h2;
    frame1[2][10] = 3'h2;
    frame1[2][11] = 3'h1;
    frame1[2][12] = 3'h1;
    frame1[2][13] = 3'h0;
    frame1[2][14] = 3'h0;
    frame1[2][15] = 3'h0;
    frame1[2][16] = 3'h0;
    frame1[2][17] = 3'h0;
    frame1[2][18] = 3'h0;
    frame1[2][19] = 3'h0;
    frame1[2][20] = 3'h0;
    frame1[2][21] = 3'h0;
    frame1[2][22] = 3'h0;
    frame1[2][23] = 3'h0;
    frame1[2][24] = 3'h0;
    // frame1[2][25] = 3'h0;
    // frame1[2][26] = 3'h0;
    // frame1[2][27] = 3'h0;
    // frame1[2][28] = 3'h0;
    // frame1[2][29] = 3'h0;
    // frame1[2][30] = 3'h0;
    // frame1[2][31] = 3'h0;
    frame1[3][0] = 3'h0;
    frame1[3][1] = 3'h0;
    frame1[3][2] = 3'h0;
    frame1[3][3] = 3'h0;
    frame1[3][4] = 3'h1;
    frame1[3][5] = 3'h1;
    frame1[3][6] = 3'h2;
    frame1[3][7] = 3'h2;
    frame1[3][8] = 3'h2;
    frame1[3][9] = 3'h2;
    frame1[3][10] = 3'h2;
    frame1[3][11] = 3'h2;
    frame1[3][12] = 3'h1;
    frame1[3][13] = 3'h0;
    frame1[3][14] = 3'h0;
    frame1[3][15] = 3'h0;
    frame1[3][16] = 3'h0;
    frame1[3][17] = 3'h0;
    frame1[3][18] = 3'h0;
    frame1[3][19] = 3'h0;
    frame1[3][20] = 3'h0;
    frame1[3][21] = 3'h0;
    frame1[3][22] = 3'h0;
    frame1[3][23] = 3'h0;
    frame1[3][24] = 3'h0;
    // frame1[3][25] = 3'h0;
    // frame1[3][26] = 3'h0;
    // frame1[3][27] = 3'h0;
    // frame1[3][28] = 3'h0;
    // frame1[3][29] = 3'h0;
    // frame1[3][30] = 3'h0;
    // frame1[3][31] = 3'h0;
    frame1[4][0] = 3'h0;
    frame1[4][1] = 3'h0;
    frame1[4][2] = 3'h0;
    frame1[4][3] = 3'h0;
    frame1[4][4] = 3'h1;
    frame1[4][5] = 3'h2;
    frame1[4][6] = 3'h2;
    frame1[4][7] = 3'h1;
    frame1[4][8] = 3'h1;
    frame1[4][9] = 3'h2;
    frame1[4][10] = 3'h2;
    frame1[4][11] = 3'h2;
    frame1[4][12] = 3'h1;
    frame1[4][13] = 3'h0;
    frame1[4][14] = 3'h0;
    frame1[4][15] = 3'h0;
    frame1[4][16] = 3'h0;
    frame1[4][17] = 3'h0;
    frame1[4][18] = 3'h0;
    frame1[4][19] = 3'h0;
    frame1[4][20] = 3'h0;
    frame1[4][21] = 3'h0;
    frame1[4][22] = 3'h0;
    frame1[4][23] = 3'h0;
    frame1[4][24] = 3'h0;
    // frame1[4][25] = 3'h0;
    // frame1[4][26] = 3'h0;
    // frame1[4][27] = 3'h0;
    // frame1[4][28] = 3'h0;
    // frame1[4][29] = 3'h0;
    // frame1[4][30] = 3'h0;
    // frame1[4][31] = 3'h0;
    frame1[5][0] = 3'h0;
    frame1[5][1] = 3'h0;
    frame1[5][2] = 3'h0;
    frame1[5][3] = 3'h0;
    frame1[5][4] = 3'h1;
    frame1[5][5] = 3'h2;
    frame1[5][6] = 3'h2;
    frame1[5][7] = 3'h1;
    frame1[5][8] = 3'h2;
    frame1[5][9] = 3'h2;
    frame1[5][10] = 3'h2;
    frame1[5][11] = 3'h2;
    frame1[5][12] = 3'h1;
    frame1[5][13] = 3'h0;
    frame1[5][14] = 3'h0;
    frame1[5][15] = 3'h0;
    frame1[5][16] = 3'h0;
    frame1[5][17] = 3'h0;
    frame1[5][18] = 3'h0;
    frame1[5][19] = 3'h0;
    frame1[5][20] = 3'h0;
    frame1[5][21] = 3'h0;
    frame1[5][22] = 3'h0;
    frame1[5][23] = 3'h0;
    frame1[5][24] = 3'h0;
    // frame1[5][25] = 3'h0;
    // frame1[5][26] = 3'h0;
    // frame1[5][27] = 3'h0;
    // frame1[5][28] = 3'h0;
    // frame1[5][29] = 3'h0;
    // frame1[5][30] = 3'h0;
    // frame1[5][31] = 3'h0;
    frame1[6][0] = 3'h0;
    frame1[6][1] = 3'h1;
    frame1[6][2] = 3'h1;
    frame1[6][3] = 3'h1;
    frame1[6][4] = 3'h1;
    frame1[6][5] = 3'h2;
    frame1[6][6] = 3'h2;
    frame1[6][7] = 3'h2;
    frame1[6][8] = 3'h2;
    frame1[6][9] = 3'h2;
    frame1[6][10] = 3'h2;
    frame1[6][11] = 3'h3;
    frame1[6][12] = 3'h1;
    frame1[6][13] = 3'h0;
    frame1[6][14] = 3'h0;
    frame1[6][15] = 3'h0;
    frame1[6][16] = 3'h0;
    frame1[6][17] = 3'h0;
    frame1[6][18] = 3'h0;
    frame1[6][19] = 3'h0;
    frame1[6][20] = 3'h0;
    frame1[6][21] = 3'h0;
    frame1[6][22] = 3'h0;
    frame1[6][23] = 3'h0;
    frame1[6][24] = 3'h0;
    // frame1[6][25] = 3'h0;
    // frame1[6][26] = 3'h0;
    // frame1[6][27] = 3'h0;
    // frame1[6][28] = 3'h0;
    // frame1[6][29] = 3'h0;
    // frame1[6][30] = 3'h0;
    // frame1[6][31] = 3'h0;
    frame1[7][0] = 3'h0;
    frame1[7][1] = 3'h1;
    frame1[7][2] = 3'h1;
    frame1[7][3] = 3'h1;
    frame1[7][4] = 3'h1;
    frame1[7][5] = 3'h1;
    frame1[7][6] = 3'h2;
    frame1[7][7] = 3'h2;
    frame1[7][8] = 3'h2;
    frame1[7][9] = 3'h2;
    frame1[7][10] = 3'h3;
    frame1[7][11] = 3'h3;
    frame1[7][12] = 3'h1;
    frame1[7][13] = 3'h0;
    frame1[7][14] = 3'h0;
    frame1[7][15] = 3'h0;
    frame1[7][16] = 3'h0;
    frame1[7][17] = 3'h0;
    frame1[7][18] = 3'h0;
    frame1[7][19] = 3'h0;
    frame1[7][20] = 3'h0;
    frame1[7][21] = 3'h0;
    frame1[7][22] = 3'h0;
    frame1[7][23] = 3'h0;
    frame1[7][24] = 3'h0;
    // frame1[7][25] = 3'h0;
    // frame1[7][26] = 3'h0;
    // frame1[7][27] = 3'h0;
    // frame1[7][28] = 3'h0;
    // frame1[7][29] = 3'h0;
    // frame1[7][30] = 3'h0;
    // frame1[7][31] = 3'h0;
    frame1[8][0] = 3'h0;
    frame1[8][1] = 3'h0;
    frame1[8][2] = 3'h0;
    frame1[8][3] = 3'h0;
    frame1[8][4] = 3'h0;
    frame1[8][5] = 3'h0;
    frame1[8][6] = 3'h1;
    frame1[8][7] = 3'h1;
    frame1[8][8] = 3'h1;
    frame1[8][9] = 3'h3;
    frame1[8][10] = 3'h3;
    frame1[8][11] = 3'h2;
    frame1[8][12] = 3'h1;
    frame1[8][13] = 3'h0;
    frame1[8][14] = 3'h0;
    frame1[8][15] = 3'h0;
    frame1[8][16] = 3'h0;
    frame1[8][17] = 3'h0;
    frame1[8][18] = 3'h0;
    frame1[8][19] = 3'h0;
    frame1[8][20] = 3'h0;
    frame1[8][21] = 3'h0;
    frame1[8][22] = 3'h0;
    frame1[8][23] = 3'h0;
    frame1[8][24] = 3'h0;
    // frame1[8][25] = 3'h0;
    // frame1[8][26] = 3'h0;
    // frame1[8][27] = 3'h0;
    // frame1[8][28] = 3'h0;
    // frame1[8][29] = 3'h0;
    // frame1[8][30] = 3'h0;
    // frame1[8][31] = 3'h0;
    frame1[9][0] = 3'h0;
    frame1[9][1] = 3'h0;
    frame1[9][2] = 3'h0;
    frame1[9][3] = 3'h0;
    frame1[9][4] = 3'h0;
    frame1[9][5] = 3'h0;
    frame1[9][6] = 3'h0;
    frame1[9][7] = 3'h0;
    frame1[9][8] = 3'h1;
    frame1[9][9] = 3'h3;
    frame1[9][10] = 3'h2;
    frame1[9][11] = 3'h2;
    frame1[9][12] = 3'h1;
    frame1[9][13] = 3'h0;
    frame1[9][14] = 3'h0;
    frame1[9][15] = 3'h0;
    frame1[9][16] = 3'h0;
    frame1[9][17] = 3'h0;
    frame1[9][18] = 3'h0;
    frame1[9][19] = 3'h0;
    frame1[9][20] = 3'h0;
    frame1[9][21] = 3'h0;
    frame1[9][22] = 3'h0;
    frame1[9][23] = 3'h0;
    frame1[9][24] = 3'h0;
    // frame1[9][25] = 3'h0;
    // frame1[9][26] = 3'h0;
    // frame1[9][27] = 3'h0;
    // frame1[9][28] = 3'h0;
    // frame1[9][29] = 3'h0;
    // frame1[9][30] = 3'h0;
    // frame1[9][31] = 3'h0;
    frame1[10][0] = 3'h0;
    frame1[10][1] = 3'h0;
    frame1[10][2] = 3'h0;
    frame1[10][3] = 3'h0;
    frame1[10][4] = 3'h0;
    frame1[10][5] = 3'h0;
    frame1[10][6] = 3'h0;
    frame1[10][7] = 3'h0;
    frame1[10][8] = 3'h1;
    frame1[10][9] = 3'h2;
    frame1[10][10] = 3'h2;
    frame1[10][11] = 3'h2;
    frame1[10][12] = 3'h1;
    frame1[10][13] = 3'h0;
    frame1[10][14] = 3'h0;
    frame1[10][15] = 3'h0;
    frame1[10][16] = 3'h0;
    frame1[10][17] = 3'h0;
    frame1[10][18] = 3'h0;
    frame1[10][19] = 3'h0;
    frame1[10][20] = 3'h0;
    frame1[10][21] = 3'h0;
    frame1[10][22] = 3'h0;
    frame1[10][23] = 3'h0;
    frame1[10][24] = 3'h0;
    // frame1[10][25] = 3'h0;
    // frame1[10][26] = 3'h0;
    // frame1[10][27] = 3'h0;
    // frame1[10][28] = 3'h0;
    // frame1[10][29] = 3'h0;
    // frame1[10][30] = 3'h0;
    // frame1[10][31] = 3'h0;
    frame1[11][0] = 3'h0;
    frame1[11][1] = 3'h0;
    frame1[11][2] = 3'h0;
    frame1[11][3] = 3'h0;
    frame1[11][4] = 3'h0;
    frame1[11][5] = 3'h0;
    frame1[11][6] = 3'h0;
    frame1[11][7] = 3'h0;
    frame1[11][8] = 3'h1;
    frame1[11][9] = 3'h2;
    frame1[11][10] = 3'h2;
    frame1[11][11] = 3'h2;
    frame1[11][12] = 3'h1;
    frame1[11][13] = 3'h0;
    frame1[11][14] = 3'h0;
    frame1[11][15] = 3'h0;
    frame1[11][16] = 3'h0;
    frame1[11][17] = 3'h0;
    frame1[11][18] = 3'h0;
    frame1[11][19] = 3'h0;
    frame1[11][20] = 3'h0;
    frame1[11][21] = 3'h0;
    frame1[11][22] = 3'h0;
    frame1[11][23] = 3'h0;
    frame1[11][24] = 3'h0;
    // frame1[11][25] = 3'h0;
    // frame1[11][26] = 3'h0;
    // frame1[11][27] = 3'h0;
    // frame1[11][28] = 3'h0;
    // frame1[11][29] = 3'h0;
    // frame1[11][30] = 3'h0;
    // frame1[11][31] = 3'h0;
    frame1[12][0] = 3'h0;
    frame1[12][1] = 3'h0;
    frame1[12][2] = 3'h0;
    frame1[12][3] = 3'h0;
    frame1[12][4] = 3'h0;
    frame1[12][5] = 3'h0;
    frame1[12][6] = 3'h0;
    frame1[12][7] = 3'h0;
    frame1[12][8] = 3'h1;
    frame1[12][9] = 3'h2;
    frame1[12][10] = 3'h2;
    frame1[12][11] = 3'h2;
    frame1[12][12] = 3'h1;
    frame1[12][13] = 3'h0;
    frame1[12][14] = 3'h0;
    frame1[12][15] = 3'h0;
    frame1[12][16] = 3'h0;
    frame1[12][17] = 3'h0;
    frame1[12][18] = 3'h0;
    frame1[12][19] = 3'h0;
    frame1[12][20] = 3'h0;
    frame1[12][21] = 3'h0;
    frame1[12][22] = 3'h0;
    frame1[12][23] = 3'h0;
    frame1[12][24] = 3'h0;
    // frame1[12][25] = 3'h0;
    // frame1[12][26] = 3'h0;
    // frame1[12][27] = 3'h0;
    // frame1[12][28] = 3'h0;
    // frame1[12][29] = 3'h0;
    // frame1[12][30] = 3'h0;
    // frame1[12][31] = 3'h0;
    frame1[13][0] = 3'h0;
    frame1[13][1] = 3'h0;
    frame1[13][2] = 3'h0;
    frame1[13][3] = 3'h0;
    frame1[13][4] = 3'h0;
    frame1[13][5] = 3'h0;
    frame1[13][6] = 3'h0;
    frame1[13][7] = 3'h0;
    frame1[13][8] = 3'h1;
    frame1[13][9] = 3'h2;
    frame1[13][10] = 3'h2;
    frame1[13][11] = 3'h2;
    frame1[13][12] = 3'h1;
    frame1[13][13] = 3'h0;
    frame1[13][14] = 3'h0;
    frame1[13][15] = 3'h0;
    frame1[13][16] = 3'h0;
    frame1[13][17] = 3'h0;
    frame1[13][18] = 3'h0;
    frame1[13][19] = 3'h0;
    frame1[13][20] = 3'h0;
    frame1[13][21] = 3'h0;
    frame1[13][22] = 3'h0;
    frame1[13][23] = 3'h0;
    frame1[13][24] = 3'h0;
    // frame1[13][25] = 3'h0;
    // frame1[13][26] = 3'h0;
    // frame1[13][27] = 3'h0;
    // frame1[13][28] = 3'h0;
    // frame1[13][29] = 3'h0;
    // frame1[13][30] = 3'h0;
    // frame1[13][31] = 3'h0;
    frame1[14][0] = 3'h0;
    frame1[14][1] = 3'h0;
    frame1[14][2] = 3'h0;
    frame1[14][3] = 3'h0;
    frame1[14][4] = 3'h0;
    frame1[14][5] = 3'h0;
    frame1[14][6] = 3'h0;
    frame1[14][7] = 3'h1;
    frame1[14][8] = 3'h1;
    frame1[14][9] = 3'h2;
    frame1[14][10] = 3'h2;
    frame1[14][11] = 3'h2;
    frame1[14][12] = 3'h1;
    frame1[14][13] = 3'h1;
    frame1[14][14] = 3'h0;
    frame1[14][15] = 3'h0;
    frame1[14][16] = 3'h0;
    frame1[14][17] = 3'h0;
    frame1[14][18] = 3'h0;
    frame1[14][19] = 3'h0;
    frame1[14][20] = 3'h0;
    frame1[14][21] = 3'h0;
    frame1[14][22] = 3'h0;
    frame1[14][23] = 3'h0;
    frame1[14][24] = 3'h0;
    // frame1[14][25] = 3'h0;
    // frame1[14][26] = 3'h0;
    // frame1[14][27] = 3'h0;
    // frame1[14][28] = 3'h0;
    // frame1[14][29] = 3'h0;
    // frame1[14][30] = 3'h0;
    // frame1[14][31] = 3'h0;
    frame1[15][0] = 3'h0;
    frame1[15][1] = 3'h0;
    frame1[15][2] = 3'h0;
    frame1[15][3] = 3'h0;
    frame1[15][4] = 3'h0;
    frame1[15][5] = 3'h0;
    frame1[15][6] = 3'h1;
    frame1[15][7] = 3'h1;
    frame1[15][8] = 3'h4;
    frame1[15][9] = 3'h4;
    frame1[15][10] = 3'h4;
    frame1[15][11] = 3'h2;
    frame1[15][12] = 3'h2;
    frame1[15][13] = 3'h1;
    frame1[15][14] = 3'h1;
    frame1[15][15] = 3'h1;
    frame1[15][16] = 3'h1;
    frame1[15][17] = 3'h1;
    frame1[15][18] = 3'h1;
    frame1[15][19] = 3'h1;
    frame1[15][20] = 3'h0;
    frame1[15][21] = 3'h0;
    frame1[15][22] = 3'h0;
    frame1[15][23] = 3'h0;
    frame1[15][24] = 3'h0;
    // frame1[15][25] = 3'h0;
    // frame1[15][26] = 3'h0;
    // frame1[15][27] = 3'h0;
    // frame1[15][28] = 3'h1;
    // frame1[15][29] = 3'h1;
    // frame1[15][30] = 3'h1;
    // frame1[15][31] = 3'h0;
    frame1[16][0] = 3'h0;
    frame1[16][1] = 3'h0;
    frame1[16][2] = 3'h0;
    frame1[16][3] = 3'h0;
    frame1[16][4] = 3'h0;
    frame1[16][5] = 3'h1;
    frame1[16][6] = 3'h1;
    frame1[16][7] = 3'h4;
    frame1[16][8] = 3'h4;
    frame1[16][9] = 3'h4;
    frame1[16][10] = 3'h5;
    frame1[16][11] = 3'h5;
    frame1[16][12] = 3'h5;
    frame1[16][13] = 3'h5;
    frame1[16][14] = 3'h5;
    frame1[16][15] = 3'h5;
    frame1[16][16] = 3'h5;
    frame1[16][17] = 3'h5;
    frame1[16][18] = 3'h5;
    frame1[16][19] = 3'h1;
    frame1[16][20] = 3'h1;
    frame1[16][21] = 3'h1;
    frame1[16][22] = 3'h1;
    frame1[16][23] = 3'h1;
    frame1[16][24] = 3'h0;
    // frame1[16][25] = 3'h0;
    // frame1[16][26] = 3'h1;
    // frame1[16][27] = 3'h1;
    // frame1[16][28] = 3'h1;
    // frame1[16][29] = 3'h5;
    // frame1[16][30] = 3'h1;
    // frame1[16][31] = 3'h0;
    frame1[17][0] = 3'h0;
    frame1[17][1] = 3'h0;
    frame1[17][2] = 3'h0;
    frame1[17][3] = 3'h0;
    frame1[17][4] = 3'h1;
    frame1[17][5] = 3'h1;
    frame1[17][6] = 3'h4;
    frame1[17][7] = 3'h4;
    frame1[17][8] = 3'h4;
    frame1[17][9] = 3'h5;
    frame1[17][10] = 3'h5;
    frame1[17][11] = 3'h5;
    frame1[17][12] = 3'h5;
    frame1[17][13] = 3'h5;
    frame1[17][14] = 3'h5;
    frame1[17][15] = 3'h5;
    frame1[17][16] = 3'h5;
    frame1[17][17] = 3'h5;
    frame1[17][18] = 3'h5;
    frame1[17][19] = 3'h5;
    frame1[17][20] = 3'h5;
    frame1[17][21] = 3'h5;
    frame1[17][22] = 3'h5;
    frame1[17][23] = 3'h1;
    frame1[17][24] = 3'h1;
    // frame1[17][25] = 3'h1;
    // frame1[17][26] = 3'h1;
    // frame1[17][27] = 3'h5;
    // frame1[17][28] = 3'h5;
    // frame1[17][29] = 3'h5;
    // frame1[17][30] = 3'h1;
    // frame1[17][31] = 3'h0;
    frame1[18][0] = 3'h0;
    frame1[18][1] = 3'h0;
    frame1[18][2] = 3'h0;
    frame1[18][3] = 3'h0;
    frame1[18][4] = 3'h1;
    frame1[18][5] = 3'h4;
    frame1[18][6] = 3'h4;
    frame1[18][7] = 3'h4;
    frame1[18][8] = 3'h5;
    frame1[18][9] = 3'h5;
    frame1[18][10] = 3'h5;
    frame1[18][11] = 3'h5;
    frame1[18][12] = 3'h5;
    frame1[18][13] = 3'h2;
    frame1[18][14] = 3'h2;
    frame1[18][15] = 3'h5;
    frame1[18][16] = 3'h5;
    frame1[18][17] = 3'h5;
    frame1[18][18] = 3'h5;
    frame1[18][19] = 3'h5;
    frame1[18][20] = 3'h5;
    frame1[18][21] = 3'h5;
    frame1[18][22] = 3'h5;
    frame1[18][23] = 3'h5;
    frame1[18][24] = 3'h5;
    // frame1[18][25] = 3'h5;
    // frame1[18][26] = 3'h5;
    // frame1[18][27] = 3'h5;
    // frame1[18][28] = 3'h5;
    // frame1[18][29] = 3'h5;
    // frame1[18][30] = 3'h1;
    // frame1[18][31] = 3'h0;
    frame1[19][0] = 3'h0;
    frame1[19][1] = 3'h0;
    frame1[19][2] = 3'h0;
    frame1[19][3] = 3'h0;
    frame1[19][4] = 3'h1;
    frame1[19][5] = 3'h4;
    frame1[19][6] = 3'h4;
    frame1[19][7] = 3'h4;
    frame1[19][8] = 3'h5;
    frame1[19][9] = 3'h5;
    frame1[19][10] = 3'h5;
    frame1[19][11] = 3'h5;
    frame1[19][12] = 3'h5;
    frame1[19][13] = 3'h1;
    frame1[19][14] = 3'h2;
    frame1[19][15] = 3'h2;
    frame1[19][16] = 3'h5;
    frame1[19][17] = 3'h5;
    frame1[19][18] = 3'h5;
    frame1[19][19] = 3'h5;
    frame1[19][20] = 3'h5;
    frame1[19][21] = 3'h5;
    frame1[19][22] = 3'h5;
    frame1[19][23] = 3'h5;
    frame1[19][24] = 3'h5;
    // frame1[19][25] = 3'h5;
    // frame1[19][26] = 3'h5;
    // frame1[19][27] = 3'h5;
    // frame1[19][28] = 3'h5;
    // frame1[19][29] = 3'h1;
    // frame1[19][30] = 3'h1;
    // frame1[19][31] = 3'h0;
    frame1[20][0] = 3'h0;
    frame1[20][1] = 3'h0;
    frame1[20][2] = 3'h0;
    frame1[20][3] = 3'h0;
    frame1[20][4] = 3'h1;
    frame1[20][5] = 3'h4;
    frame1[20][6] = 3'h4;
    frame1[20][7] = 3'h4;
    frame1[20][8] = 3'h4;
    frame1[20][9] = 3'h5;
    frame1[20][10] = 3'h5;
    frame1[20][11] = 3'h5;
    frame1[20][12] = 3'h5;
    frame1[20][13] = 3'h5;
    frame1[20][14] = 3'h5;
    frame1[20][15] = 3'h5;
    frame1[20][16] = 3'h1;
    frame1[20][17] = 3'h2;
    frame1[20][18] = 3'h2;
    frame1[20][19] = 3'h2;
    frame1[20][20] = 3'h2;
    frame1[20][21] = 3'h2;
    frame1[20][22] = 3'h2;
    frame1[20][23] = 3'h2;
    frame1[20][24] = 3'h2;
    // frame1[20][25] = 3'h1;
    // frame1[20][26] = 3'h3;
    // frame1[20][27] = 3'h1;
    // frame1[20][28] = 3'h1;
    // frame1[20][29] = 3'h0;
    // frame1[20][30] = 3'h0;
    // frame1[20][31] = 3'h0;
    frame1[21][0] = 3'h0;
    frame1[21][1] = 3'h0;
    frame1[21][2] = 3'h0;
    frame1[21][3] = 3'h0;
    frame1[21][4] = 3'h1;
    frame1[21][5] = 3'h1;
    frame1[21][6] = 3'h1;
    frame1[21][7] = 3'h4;
    frame1[21][8] = 3'h4;
    frame1[21][9] = 3'h4;
    frame1[21][10] = 3'h5;
    frame1[21][11] = 3'h5;
    frame1[21][12] = 3'h5;
    frame1[21][13] = 3'h5;
    frame1[21][14] = 3'h5;
    frame1[21][15] = 3'h5;
    frame1[21][16] = 3'h5;
    frame1[21][17] = 3'h1;
    frame1[21][18] = 3'h1;
    frame1[21][19] = 3'h1;
    frame1[21][20] = 3'h1;
    frame1[21][21] = 3'h1;
    frame1[21][22] = 3'h1;
    frame1[21][23] = 3'h1;
    frame1[21][24] = 3'h3;
    // frame1[21][25] = 3'h1;
    // frame1[21][26] = 3'h1;
    // frame1[21][27] = 3'h0;
    // frame1[21][28] = 3'h0;
    // frame1[21][29] = 3'h0;
    // frame1[21][30] = 3'h0;
    // frame1[21][31] = 3'h0;
    frame1[22][0] = 3'h0;
    frame1[22][1] = 3'h0;
    frame1[22][2] = 3'h0;
    frame1[22][3] = 3'h0;
    frame1[22][4] = 3'h0;
    frame1[22][5] = 3'h0;
    frame1[22][6] = 3'h1;
    frame1[22][7] = 3'h1;
    frame1[22][8] = 3'h4;
    frame1[22][9] = 3'h4;
    frame1[22][10] = 3'h4;
    frame1[22][11] = 3'h5;
    frame1[22][12] = 3'h5;
    frame1[22][13] = 3'h5;
    frame1[22][14] = 3'h5;
    frame1[22][15] = 3'h5;
    frame1[22][16] = 3'h5;
    frame1[22][17] = 3'h3;
    frame1[22][18] = 3'h3;
    frame1[22][19] = 3'h3;
    frame1[22][20] = 3'h3;
    frame1[22][21] = 3'h3;
    frame1[22][22] = 3'h3;
    frame1[22][23] = 3'h3;
    frame1[22][24] = 3'h1;
    // frame1[22][25] = 3'h1;
    // frame1[22][26] = 3'h0;
    // frame1[22][27] = 3'h0;
    // frame1[22][28] = 3'h0;
    // frame1[22][29] = 3'h0;
    // frame1[22][30] = 3'h0;
    // frame1[22][31] = 3'h0;
    frame1[23][0] = 3'h0;
    frame1[23][1] = 3'h0;
    frame1[23][2] = 3'h0;
    frame1[23][3] = 3'h0;
    frame1[23][4] = 3'h0;
    frame1[23][5] = 3'h0;
    frame1[23][6] = 3'h0;
    frame1[23][7] = 3'h1;
    frame1[23][8] = 3'h1;
    frame1[23][9] = 3'h4;
    frame1[23][10] = 3'h4;
    frame1[23][11] = 3'h4;
    frame1[23][12] = 3'h4;
    frame1[23][13] = 3'h4;
    frame1[23][14] = 3'h4;
    frame1[23][15] = 3'h4;
    frame1[23][16] = 3'h4;
    frame1[23][17] = 3'h4;
    frame1[23][18] = 3'h4;
    frame1[23][19] = 3'h4;
    frame1[23][20] = 3'h4;
    frame1[23][21] = 3'h4;
    frame1[23][22] = 3'h1;
    frame1[23][23] = 3'h1;
    frame1[23][24] = 3'h1;
    // frame1[23][25] = 3'h0;
    // frame1[23][26] = 3'h0;
    // frame1[23][27] = 3'h0;
    // frame1[23][28] = 3'h0;
    // frame1[23][29] = 3'h0;
    // frame1[23][30] = 3'h0;
    // frame1[23][31] = 3'h0;
    frame1[24][0] = 3'h0;
    frame1[24][1] = 3'h0;
    frame1[24][2] = 3'h0;
    frame1[24][3] = 3'h0;
    frame1[24][4] = 3'h0;
    frame1[24][5] = 3'h0;
    frame1[24][6] = 3'h0;
    frame1[24][7] = 3'h0;
    frame1[24][8] = 3'h1;
    frame1[24][9] = 3'h1;
    frame1[24][10] = 3'h1;
    frame1[24][11] = 3'h1;
    frame1[24][12] = 3'h5;
    frame1[24][13] = 3'h5;
    frame1[24][14] = 3'h5;
    frame1[24][15] = 3'h1;
    frame1[24][16] = 3'h1;
    frame1[24][17] = 3'h1;
    frame1[24][18] = 3'h1;
    frame1[24][19] = 3'h1;
    frame1[24][20] = 3'h1;
    frame1[24][21] = 3'h1;
    frame1[24][22] = 3'h0;
    frame1[24][23] = 3'h0;
    frame1[24][24] = 3'h0;
    // frame1[24][25] = 3'h0;
    // frame1[24][26] = 3'h0;
    // frame1[24][27] = 3'h0;
    // frame1[24][28] = 3'h0;
    // frame1[24][29] = 3'h0;
    // frame1[24][30] = 3'h0;
    // frame1[24][31] = 3'h0;
    // frame1[25][0] = 3'h0;
    // frame1[25][1] = 3'h0;
    // frame1[25][2] = 3'h0;
    // frame1[25][3] = 3'h0;
    // frame1[25][4] = 3'h0;
    // frame1[25][5] = 3'h0;
    // frame1[25][6] = 3'h0;
    // frame1[25][7] = 3'h0;
    // frame1[25][8] = 3'h0;
    // frame1[25][9] = 3'h0;
    // frame1[25][10] = 3'h1;
    // frame1[25][11] = 3'h1;
    // frame1[25][12] = 3'h1;
    // frame1[25][13] = 3'h1;
    // frame1[25][14] = 3'h1;
    // frame1[25][15] = 3'h1;
    // frame1[25][16] = 3'h0;
    // frame1[25][17] = 3'h1;
    // frame1[25][18] = 3'h0;
    // frame1[25][19] = 3'h0;
    // frame1[25][20] = 3'h0;
    // frame1[25][21] = 3'h0;
    // frame1[25][22] = 3'h0;
    // frame1[25][23] = 3'h0;
    // frame1[25][24] = 3'h0;
    // frame1[25][25] = 3'h0;
    // frame1[25][26] = 3'h0;
    // frame1[25][27] = 3'h0;
    // frame1[25][28] = 3'h0;
    // frame1[25][29] = 3'h0;
    // frame1[25][30] = 3'h0;
    // frame1[25][31] = 3'h0;
    // frame1[26][0] = 3'h0;
    // frame1[26][1] = 3'h0;
    // frame1[26][2] = 3'h0;
    // frame1[26][3] = 3'h0;
    // frame1[26][4] = 3'h0;
    // frame1[26][5] = 3'h0;
    // frame1[26][6] = 3'h0;
    // frame1[26][7] = 3'h0;
    // frame1[26][8] = 3'h0;
    // frame1[26][9] = 3'h0;
    // frame1[26][10] = 3'h0;
    // frame1[26][11] = 3'h0;
    // frame1[26][12] = 3'h0;
    // frame1[26][13] = 3'h1;
    // frame1[26][14] = 3'h0;
    // frame1[26][15] = 3'h0;
    // frame1[26][16] = 3'h0;
    // frame1[26][17] = 3'h1;
    // frame1[26][18] = 3'h0;
    // frame1[26][19] = 3'h0;
    // frame1[26][20] = 3'h0;
    // frame1[26][21] = 3'h0;
    // frame1[26][22] = 3'h0;
    // frame1[26][23] = 3'h0;
    // frame1[26][24] = 3'h0;
    // frame1[26][25] = 3'h0;
    // frame1[26][26] = 3'h0;
    // frame1[26][27] = 3'h0;
    // frame1[26][28] = 3'h0;
    // frame1[26][29] = 3'h0;
    // frame1[26][30] = 3'h0;
    // frame1[26][31] = 3'h0;
    // frame1[27][0] = 3'h0;
    // frame1[27][1] = 3'h0;
    // frame1[27][2] = 3'h0;
    // frame1[27][3] = 3'h0;
    // frame1[27][4] = 3'h0;
    // frame1[27][5] = 3'h0;
    // frame1[27][6] = 3'h0;
    // frame1[27][7] = 3'h0;
    // frame1[27][8] = 3'h0;
    // frame1[27][9] = 3'h0;
    // frame1[27][10] = 3'h0;
    // frame1[27][11] = 3'h0;
    // frame1[27][12] = 3'h0;
    // frame1[27][13] = 3'h1;
    // frame1[27][14] = 3'h0;
    // frame1[27][15] = 3'h0;
    // frame1[27][16] = 3'h0;
    // frame1[27][17] = 3'h1;
    // frame1[27][18] = 3'h0;
    // frame1[27][19] = 3'h0;
    // frame1[27][20] = 3'h0;
    // frame1[27][21] = 3'h0;
    // frame1[27][22] = 3'h0;
    // frame1[27][23] = 3'h0;
    // frame1[27][24] = 3'h0;
    // frame1[27][25] = 3'h0;
    // frame1[27][26] = 3'h0;
    // frame1[27][27] = 3'h0;
    // frame1[27][28] = 3'h0;
    // frame1[27][29] = 3'h0;
    // frame1[27][30] = 3'h0;
    // frame1[27][31] = 3'h0;
    // frame1[28][0] = 3'h0;
    // frame1[28][1] = 3'h0;
    // frame1[28][2] = 3'h0;
    // frame1[28][3] = 3'h0;
    // frame1[28][4] = 3'h0;
    // frame1[28][5] = 3'h0;
    // frame1[28][6] = 3'h0;
    // frame1[28][7] = 3'h0;
    // frame1[28][8] = 3'h0;
    // frame1[28][9] = 3'h0;
    // frame1[28][10] = 3'h0;
    // frame1[28][11] = 3'h0;
    // frame1[28][12] = 3'h0;
    // frame1[28][13] = 3'h1;
    // frame1[28][14] = 3'h0;
    // frame1[28][15] = 3'h0;
    // frame1[28][16] = 3'h0;
    // frame1[28][17] = 3'h1;
    // frame1[28][18] = 3'h0;
    // frame1[28][19] = 3'h0;
    // frame1[28][20] = 3'h0;
    // frame1[28][21] = 3'h0;
    // frame1[28][22] = 3'h0;
    // frame1[28][23] = 3'h0;
    // frame1[28][24] = 3'h0;
    // frame1[28][25] = 3'h0;
    // frame1[28][26] = 3'h0;
    // frame1[28][27] = 3'h0;
    // frame1[28][28] = 3'h0;
    // frame1[28][29] = 3'h0;
    // frame1[28][30] = 3'h0;
    // frame1[28][31] = 3'h0;
    // frame1[29][0] = 3'h0;
    // frame1[29][1] = 3'h0;
    // frame1[29][2] = 3'h0;
    // frame1[29][3] = 3'h0;
    // frame1[29][4] = 3'h0;
    // frame1[29][5] = 3'h0;
    // frame1[29][6] = 3'h0;
    // frame1[29][7] = 3'h0;
    // frame1[29][8] = 3'h0;
    // frame1[29][9] = 3'h0;
    // frame1[29][10] = 3'h0;
    // frame1[29][11] = 3'h0;
    // frame1[29][12] = 3'h0;
    // frame1[29][13] = 3'h1;
    // frame1[29][14] = 3'h0;
    // frame1[29][15] = 3'h0;
    // frame1[29][16] = 3'h0;
    // frame1[29][17] = 3'h1;
    // frame1[29][18] = 3'h0;
    // frame1[29][19] = 3'h0;
    // frame1[29][20] = 3'h0;
    // frame1[29][21] = 3'h0;
    // frame1[29][22] = 3'h0;
    // frame1[29][23] = 3'h0;
    // frame1[29][24] = 3'h0;
    // frame1[29][25] = 3'h0;
    // frame1[29][26] = 3'h0;
    // frame1[29][27] = 3'h0;
    // frame1[29][28] = 3'h0;
    // frame1[29][29] = 3'h0;
    // frame1[29][30] = 3'h0;
    // frame1[29][31] = 3'h0;
    // frame1[30][0] = 3'h0;
    // frame1[30][1] = 3'h0;
    // frame1[30][2] = 3'h0;
    // frame1[30][3] = 3'h0;
    // frame1[30][4] = 3'h0;
    // frame1[30][5] = 3'h0;
    // frame1[30][6] = 3'h0;
    // frame1[30][7] = 3'h0;
    // frame1[30][8] = 3'h0;
    // frame1[30][9] = 3'h0;
    // frame1[30][10] = 3'h0;
    // frame1[30][11] = 3'h1;
    // frame1[30][12] = 3'h1;
    // frame1[30][13] = 3'h1;
    // frame1[30][14] = 3'h0;
    // frame1[30][15] = 3'h0;
    // frame1[30][16] = 3'h1;
    // frame1[30][17] = 3'h1;
    // frame1[30][18] = 3'h0;
    // frame1[30][19] = 3'h0;
    // frame1[30][20] = 3'h0;
    // frame1[30][21] = 3'h0;
    // frame1[30][22] = 3'h0;
    // frame1[30][23] = 3'h0;
    // frame1[30][24] = 3'h0;
    // frame1[30][25] = 3'h0;
    // frame1[30][26] = 3'h0;
    // frame1[30][27] = 3'h0;
    // frame1[30][28] = 3'h0;
    // frame1[30][29] = 3'h0;
    // frame1[30][30] = 3'h0;
    // frame1[30][31] = 3'h0;
    // frame1[31][0] = 3'h0;
    // frame1[31][1] = 3'h0;
    // frame1[31][2] = 3'h0;
    // frame1[31][3] = 3'h0;
    // frame1[31][4] = 3'h0;
    // frame1[31][5] = 3'h0;
    // frame1[31][6] = 3'h0;
    // frame1[31][7] = 3'h0;
    // frame1[31][8] = 3'h0;
    // frame1[31][9] = 3'h0;
    // frame1[31][10] = 3'h1;
    // frame1[31][11] = 3'h1;
    // frame1[31][12] = 3'h1;
    // frame1[31][13] = 3'h1;
    // frame1[31][14] = 3'h0;
    // frame1[31][15] = 3'h1;
    // frame1[31][16] = 3'h1;
    // frame1[31][17] = 3'h1;
    // frame1[31][18] = 3'h0;
    // frame1[31][19] = 3'h0;
    // frame1[31][20] = 3'h0;
    // frame1[31][21] = 3'h0;
    // frame1[31][22] = 3'h0;
    // frame1[31][23] = 3'h0;
    // frame1[31][24] = 3'h0;
    // frame1[31][25] = 3'h0;
    // frame1[31][26] = 3'h0;
    // frame1[31][27] = 3'h0;
    // frame1[31][28] = 3'h0;
    // frame1[31][29] = 3'h0;
    // frame1[31][30] = 3'h0;
    // frame1[31][31] = 3'h0;
end