reg [5:0] frame1[7:0][31:0];
initial begin
    frame1[0][0] = 6'd0;
    frame1[1][0] = 6'd0;
    frame1[2][0] = 6'd0;
    frame1[3][0] = 6'd0;
    frame1[4][0] = 6'd0;
    frame1[5][0] = 6'd0;
    frame1[6][0] = 6'd0;
    frame1[7][0] = 6'd0;
    frame1[0][1] = 6'd0;
    frame1[1][1] = 6'd0;
    frame1[2][1] = 6'd0;
    frame1[3][1] = 6'd0;
    frame1[4][1] = 6'd0;
    frame1[5][1] = 6'd0;
    frame1[6][1] = 6'd0;
    frame1[7][1] = 6'd0;
    frame1[0][2] = 6'd0;
    frame1[1][2] = 6'd3;
    frame1[2][2] = 6'd4;
    frame1[3][2] = 6'd0;
    frame1[4][2] = 6'd0;
    frame1[5][2] = 6'd0;
    frame1[6][2] = 6'd0;
    frame1[7][2] = 6'd0;
    frame1[0][3] = 6'd0;
    frame1[1][3] = 6'd7;
    frame1[2][3] = 6'd1;
    frame1[3][3] = 6'd0;
    frame1[4][3] = 6'd0;
    frame1[5][3] = 6'd0;
    frame1[6][3] = 6'd0;
    frame1[7][3] = 6'd0;
    frame1[0][4] = 6'd0;
    frame1[1][4] = 6'd13;
    frame1[2][4] = 6'd5;
    frame1[3][4] = 6'd0;
    frame1[4][4] = 6'd0;
    frame1[5][4] = 6'd0;
    frame1[6][4] = 6'd0;
    frame1[7][4] = 6'd0;
    frame1[0][5] = 6'd0;
    frame1[1][5] = 6'd13;
    frame1[2][5] = 6'd1;
    frame1[3][5] = 6'd0;
    frame1[4][5] = 6'd0;
    frame1[5][5] = 6'd0;
    frame1[6][5] = 6'd0;
    frame1[7][5] = 6'd0;
    frame1[0][6] = 6'd0;
    frame1[1][6] = 6'd5;
    frame1[2][6] = 6'd35;
    frame1[3][6] = 6'd0;
    frame1[4][6] = 6'd0;
    frame1[5][6] = 6'd0;
    frame1[6][6] = 6'd0;
    frame1[7][6] = 6'd0;
    frame1[0][7] = 6'd0;
    frame1[1][7] = 6'd7;
    frame1[2][7] = 6'd38;
    frame1[3][7] = 6'd0;
    frame1[4][7] = 6'd0;
    frame1[5][7] = 6'd0;
    frame1[6][7] = 6'd0;
    frame1[7][7] = 6'd0;
    frame1[0][8] = 6'd0;
    frame1[1][8] = 6'd0;
    frame1[2][8] = 6'd55;
    frame1[3][8] = 6'd0;
    frame1[4][8] = 6'd0;
    frame1[5][8] = 6'd0;
    frame1[6][8] = 6'd0;
    frame1[7][8] = 6'd0;
    frame1[0][9] = 6'd0;
    frame1[1][9] = 6'd0;
    frame1[2][9] = 6'd22;
    frame1[3][9] = 6'd0;
    frame1[4][9] = 6'd0;
    frame1[5][9] = 6'd0;
    frame1[6][9] = 6'd0;
    frame1[7][9] = 6'd0;
    frame1[0][10] = 6'd0;
    frame1[1][10] = 6'd0;
    frame1[2][10] = 6'd5;
    frame1[3][10] = 6'd0;
    frame1[4][10] = 6'd0;
    frame1[5][10] = 6'd0;
    frame1[6][10] = 6'd0;
    frame1[7][10] = 6'd0;
    frame1[0][11] = 6'd0;
    frame1[1][11] = 6'd0;
    frame1[2][11] = 6'd5;
    frame1[3][11] = 6'd0;
    frame1[4][11] = 6'd0;
    frame1[5][11] = 6'd0;
    frame1[6][11] = 6'd0;
    frame1[7][11] = 6'd0;
    frame1[0][12] = 6'd0;
    frame1[1][12] = 6'd0;
    frame1[2][12] = 6'd5;
    frame1[3][12] = 6'd0;
    frame1[4][12] = 6'd0;
    frame1[5][12] = 6'd0;
    frame1[6][12] = 6'd0;
    frame1[7][12] = 6'd0;
    frame1[0][13] = 6'd0;
    frame1[1][13] = 6'd0;
    frame1[2][13] = 6'd5;
    frame1[3][13] = 6'd0;
    frame1[4][13] = 6'd0;
    frame1[5][13] = 6'd0;
    frame1[6][13] = 6'd0;
    frame1[7][13] = 6'd0;
    frame1[0][14] = 6'd0;
    frame1[1][14] = 6'd0;
    frame1[2][14] = 6'd5;
    frame1[3][14] = 6'd0;
    frame1[4][14] = 6'd0;
    frame1[5][14] = 6'd0;
    frame1[6][14] = 6'd0;
    frame1[7][14] = 6'd0;
    frame1[0][15] = 6'd0;
    frame1[1][15] = 6'd0;
    frame1[2][15] = 6'd15;
    frame1[3][15] = 6'd2;
    frame1[4][15] = 6'd0;
    frame1[5][15] = 6'd0;
    frame1[6][15] = 6'd0;
    frame1[7][15] = 6'd0;
    frame1[0][16] = 6'd0;
    frame1[1][16] = 6'd16;
    frame1[2][16] = 6'd12;
    frame1[3][16] = 6'd1;
    frame1[4][16] = 6'd4;
    frame1[5][16] = 6'd0;
    frame1[6][16] = 6'd0;
    frame1[7][16] = 6'd37;
    frame1[0][17] = 6'd0;
    frame1[1][17] = 6'd26;
    frame1[2][17] = 6'd31;
    frame1[3][17] = 6'd1;
    frame1[4][17] = 6'd1;
    frame1[5][17] = 6'd4;
    frame1[6][17] = 6'd3;
    frame1[7][17] = 6'd8;
    frame1[0][18] = 6'd0;
    frame1[1][18] = 6'd9;
    frame1[2][18] = 6'd1;
    frame1[3][18] = 6'd1;
    frame1[4][18] = 6'd1;
    frame1[5][18] = 6'd1;
    frame1[6][18] = 6'd1;
    frame1[7][18] = 6'd8;
    frame1[0][19] = 6'd0;
    frame1[1][19] = 6'd9;
    frame1[2][19] = 6'd1;
    frame1[3][19] = 6'd19;
    frame1[4][19] = 6'd1;
    frame1[5][19] = 6'd1;
    frame1[6][19] = 6'd1;
    frame1[7][19] = 6'd2;
    frame1[0][20] = 6'd0;
    frame1[1][20] = 6'd9;
    frame1[2][20] = 6'd1;
    frame1[3][20] = 6'd8;
    frame1[4][20] = 6'd1;
    frame1[5][20] = 6'd1;
    frame1[6][20] = 6'd18;
    frame1[7][20] = 6'd0;
    frame1[0][21] = 6'd0;
    frame1[1][21] = 6'd9;
    frame1[2][21] = 6'd31;
    frame1[3][21] = 6'd1;
    frame1[4][21] = 6'd5;
    frame1[5][21] = 6'd1;
    frame1[6][21] = 6'd47;
    frame1[7][21] = 6'd0;
    frame1[0][22] = 6'd0;
    frame1[1][22] = 6'd16;
    frame1[2][22] = 6'd12;
    frame1[3][22] = 6'd1;
    frame1[4][22] = 6'd2;
    frame1[5][22] = 6'd0;
    frame1[6][22] = 6'd27;
    frame1[7][22] = 6'd0;
    frame1[0][23] = 6'd0;
    frame1[1][23] = 6'd0;
    frame1[2][23] = 6'd15;
    frame1[3][23] = 6'd1;
    frame1[4][23] = 6'd42;
    frame1[5][23] = 6'd20;
    frame1[6][23] = 6'd52;
    frame1[7][23] = 6'd0;
    frame1[0][24] = 6'd0;
    frame1[1][24] = 6'd0;
    frame1[2][24] = 6'd9;
    frame1[3][24] = 6'd6;
    frame1[4][24] = 6'd25;
    frame1[5][24] = 6'd21;
    frame1[6][24] = 6'd0;
    frame1[7][24] = 6'd0;
    frame1[0][25] = 6'd0;
    frame1[1][25] = 6'd0;
    frame1[2][25] = 6'd16;
    frame1[3][25] = 6'd6;
    frame1[4][25] = 6'd6;
    frame1[5][25] = 6'd29;
    frame1[6][25] = 6'd0;
    frame1[7][25] = 6'd0;
    frame1[0][26] = 6'd0;
    frame1[1][26] = 6'd0;
    frame1[2][26] = 6'd0;
    frame1[3][26] = 6'd7;
    frame1[4][26] = 6'd2;
    frame1[5][26] = 6'd0;
    frame1[6][26] = 6'd0;
    frame1[7][26] = 6'd0;
    frame1[0][27] = 6'd0;
    frame1[1][27] = 6'd0;
    frame1[2][27] = 6'd0;
    frame1[3][27] = 6'd0;
    frame1[4][27] = 6'd0;
    frame1[5][27] = 6'd0;
    frame1[6][27] = 6'd0;
    frame1[7][27] = 6'd0;
    frame1[0][28] = 6'd0;
    frame1[1][28] = 6'd0;
    frame1[2][28] = 6'd0;
    frame1[3][28] = 6'd0;
    frame1[4][28] = 6'd0;
    frame1[5][28] = 6'd0;
    frame1[6][28] = 6'd0;
    frame1[7][28] = 6'd0;
    frame1[0][29] = 6'd0;
    frame1[1][29] = 6'd0;
    frame1[2][29] = 6'd0;
    frame1[3][29] = 6'd0;
    frame1[4][29] = 6'd0;
    frame1[5][29] = 6'd0;
    frame1[6][29] = 6'd0;
    frame1[7][29] = 6'd0;
    frame1[0][30] = 6'd0;
    frame1[1][30] = 6'd0;
    frame1[2][30] = 6'd0;
    frame1[3][30] = 6'd0;
    frame1[4][30] = 6'd0;
    frame1[5][30] = 6'd0;
    frame1[6][30] = 6'd0;
    frame1[7][30] = 6'd0;
    frame1[0][31] = 6'd0;
    frame1[1][31] = 6'd0;
    frame1[2][31] = 6'd0;
    frame1[3][31] = 6'd0;
    frame1[4][31] = 6'd0;
    frame1[5][31] = 6'd0;
    frame1[6][31] = 6'd0;
    frame1[7][31] = 6'd0;
end
