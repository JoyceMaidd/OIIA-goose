// 64×64 pixels, each 4 bits
reg [2:0] frame0 [0:15][0:15];

initial begin
    frame0[0][0] = 3'd0;
    frame0[0][1] = 3'd0;
    frame0[0][2] = 3'd0;
    frame0[0][3] = 3'd0;
    frame0[0][4] = 3'd0;
    frame0[0][5] = 3'd0;
    frame0[0][6] = 3'd0;
    frame0[0][7] = 3'd0;
    frame0[0][8] = 3'd0;
    frame0[0][9] = 3'd0;
    frame0[0][10] = 3'd0;
    frame0[0][11] = 3'd0;
    frame0[0][12] = 3'd0;
    frame0[0][13] = 3'd0;
    frame0[0][14] = 3'd0;
    frame0[0][15] = 3'd0;
    // frame0[0][16] = 3'd0;
    // frame0[0][17] = 3'd0;
    // frame0[0][18] = 3'd0;
    // frame0[0][19] = 3'd0;
    // frame0[0][20] = 3'd0;
    // frame0[0][21] = 3'd0;
    // frame0[0][22] = 3'd0;
    // frame0[0][23] = 3'd0;
    // frame0[0][24] = 3'd0;
    // frame0[0][25] = 3'd0;
    // frame0[0][26] = 3'd0;
    // frame0[0][27] = 3'd0;
    // frame0[0][28] = 3'd0;
    // frame0[0][29] = 3'd0;
    // frame0[0][30] = 3'd0;
    // frame0[0][31] = 3'd0;
    frame0[1][0] = 3'd0;
    frame0[1][1] = 3'd0;
    frame0[1][2] = 3'd0;
    frame0[1][3] = 3'd0;
    frame0[1][4] = 3'd0;
    frame0[1][5] = 3'd0;
    frame0[1][6] = 3'd0;
    frame0[1][7] = 3'd0;
    frame0[1][8] = 3'd0;
    frame0[1][9] = 3'd0;
    frame0[1][10] = 3'd0;
    frame0[1][11] = 3'd0;
    frame0[1][12] = 3'd0;
    frame0[1][13] = 3'd1;
    frame0[1][14] = 3'd1;
    frame0[1][15] = 3'd1;
    // frame0[1][16] = 3'd1;
    // frame0[1][17] = 3'd1;
    // frame0[1][18] = 3'd1;
    // frame0[1][19] = 3'd0;
    // frame0[1][20] = 3'd0;
    // frame0[1][21] = 3'd0;
    // frame0[1][22] = 3'd0;
    // frame0[1][23] = 3'd0;
    // frame0[1][24] = 3'd0;
    // frame0[1][25] = 3'd0;
    // frame0[1][26] = 3'd0;
    // frame0[1][27] = 3'd0;
    // frame0[1][28] = 3'd0;
    // frame0[1][29] = 3'd0;
    // frame0[1][30] = 3'd0;
    // frame0[1][31] = 3'd0;
    frame0[2][0] = 3'd0;
    frame0[2][1] = 3'd0;
    frame0[2][2] = 3'd0;
    frame0[2][3] = 3'd0;
    frame0[2][4] = 3'd0;
    frame0[2][5] = 3'd0;
    frame0[2][6] = 3'd0;
    frame0[2][7] = 3'd0;
    frame0[2][8] = 3'd0;
    frame0[2][9] = 3'd0;
    frame0[2][10] = 3'd0;
    frame0[2][11] = 3'd0;
    frame0[2][12] = 3'd1;
    frame0[2][13] = 3'd1;
    frame0[2][14] = 3'd2;
    frame0[2][15] = 3'd2;
    // frame0[2][16] = 3'd2;
    // frame0[2][17] = 3'd2;
    // frame0[2][18] = 3'd1;
    // frame0[2][19] = 3'd1;
    // frame0[2][20] = 3'd0;
    // frame0[2][21] = 3'd0;
    // frame0[2][22] = 3'd0;
    // frame0[2][23] = 3'd0;
    // frame0[2][24] = 3'd0;
    // frame0[2][25] = 3'd0;
    // frame0[2][26] = 3'd0;
    // frame0[2][27] = 3'd0;
    // frame0[2][28] = 3'd0;
    // frame0[2][29] = 3'd0;
    // frame0[2][30] = 3'd0;
    // frame0[2][31] = 3'd0;
    frame0[3][0] = 3'd0;
    frame0[3][1] = 3'd0;
    frame0[3][2] = 3'd0;
    frame0[3][3] = 3'd0;
    frame0[3][4] = 3'd0;
    frame0[3][5] = 3'd0;
    frame0[3][6] = 3'd0;
    frame0[3][7] = 3'd0;
    frame0[3][8] = 3'd0;
    frame0[3][9] = 3'd0;
    frame0[3][10] = 3'd0;
    frame0[3][11] = 3'd1;
    frame0[3][12] = 3'd2;
    frame0[3][13] = 3'd2;
    frame0[3][14] = 3'd2;
    frame0[3][15] = 3'd2;
    // frame0[3][16] = 3'd2;
    // frame0[3][17] = 3'd2;
    // frame0[3][18] = 3'd2;
    // frame0[3][19] = 3'd2;
    // frame0[3][20] = 3'd1;
    // frame0[3][21] = 3'd0;
    // frame0[3][22] = 3'd0;
    // frame0[3][23] = 3'd0;
    // frame0[3][24] = 3'd0;
    // frame0[3][25] = 3'd0;
    // frame0[3][26] = 3'd0;
    // frame0[3][27] = 3'd0;
    // frame0[3][28] = 3'd0;
    // frame0[3][29] = 3'd0;
    // frame0[3][30] = 3'd0;
    // frame0[3][31] = 3'd0;
    frame0[4][0] = 3'd0;
    frame0[4][1] = 3'd0;
    frame0[4][2] = 3'd0;
    frame0[4][3] = 3'd0;
    frame0[4][4] = 3'd0;
    frame0[4][5] = 3'd0;
    frame0[4][6] = 3'd0;
    frame0[4][7] = 3'd0;
    frame0[4][8] = 3'd0;
    frame0[4][9] = 3'd0;
    frame0[4][10] = 3'd0;
    frame0[4][11] = 3'd1;
    frame0[4][12] = 3'd1;
    frame0[4][13] = 3'd1;
    frame0[4][14] = 3'd2;
    frame0[4][15] = 3'd2;
    // frame0[4][16] = 3'd2;
    // frame0[4][17] = 3'd2;
    // frame0[4][18] = 3'd1;
    // frame0[4][19] = 3'd1;
    // frame0[4][20] = 3'd1;
    // frame0[4][21] = 3'd0;
    // frame0[4][22] = 3'd0;
    // frame0[4][23] = 3'd0;
    // frame0[4][24] = 3'd0;
    // frame0[4][25] = 3'd0;
    // frame0[4][26] = 3'd0;
    // frame0[4][27] = 3'd0;
    // frame0[4][28] = 3'd0;
    // frame0[4][29] = 3'd0;
    // frame0[4][30] = 3'd0;
    // frame0[4][31] = 3'd0;
    frame0[5][0] = 3'd0;
    frame0[5][1] = 3'd0;
    frame0[5][2] = 3'd0;
    frame0[5][3] = 3'd0;
    frame0[5][4] = 3'd0;
    frame0[5][5] = 3'd0;
    frame0[5][6] = 3'd0;
    frame0[5][7] = 3'd0;
    frame0[5][8] = 3'd0;
    frame0[5][9] = 3'd0;
    frame0[5][10] = 3'd0;
    frame0[5][11] = 3'd1;
    frame0[5][12] = 3'd3;
    frame0[5][13] = 3'd1;
    frame0[5][14] = 3'd2;
    frame0[5][15] = 3'd2;
    // frame0[5][16] = 3'd2;
    // frame0[5][17] = 3'd2;
    // frame0[5][18] = 3'd1;
    // frame0[5][19] = 3'd3;
    // frame0[5][20] = 3'd1;
    // frame0[5][21] = 3'd0;
    // frame0[5][22] = 3'd0;
    // frame0[5][23] = 3'd0;
    // frame0[5][24] = 3'd0;
    // frame0[5][25] = 3'd0;
    // frame0[5][26] = 3'd0;
    // frame0[5][27] = 3'd0;
    // frame0[5][28] = 3'd0;
    // frame0[5][29] = 3'd0;
    // frame0[5][30] = 3'd0;
    // frame0[5][31] = 3'd0;
    frame0[6][0] = 3'd0;
    frame0[6][1] = 3'd0;
    frame0[6][2] = 3'd0;
    frame0[6][3] = 3'd0;
    frame0[6][4] = 3'd0;
    frame0[6][5] = 3'd0;
    frame0[6][6] = 3'd0;
    frame0[6][7] = 3'd0;
    frame0[6][8] = 3'd0;
    frame0[6][9] = 3'd0;
    frame0[6][10] = 3'd0;
    frame0[6][11] = 3'd1;
    frame0[6][12] = 3'd1;
    frame0[6][13] = 3'd3;
    frame0[6][14] = 3'd2;
    frame0[6][15] = 3'd1;
    // frame0[6][16] = 3'd1;
    // frame0[6][17] = 3'd2;
    // frame0[6][18] = 3'd3;
    // frame0[6][19] = 3'd1;
    // frame0[6][20] = 3'd1;
    // frame0[6][21] = 3'd0;
    // frame0[6][22] = 3'd0;
    // frame0[6][23] = 3'd0;
    // frame0[6][24] = 3'd0;
    // frame0[6][25] = 3'd0;
    // frame0[6][26] = 3'd0;
    // frame0[6][27] = 3'd0;
    // frame0[6][28] = 3'd0;
    // frame0[6][29] = 3'd0;
    // frame0[6][30] = 3'd0;
    // frame0[6][31] = 3'd0;
    frame0[7][0] = 3'd0;
    frame0[7][1] = 3'd0;
    frame0[7][2] = 3'd0;
    frame0[7][3] = 3'd0;
    frame0[7][4] = 3'd0;
    frame0[7][5] = 3'd0;
    frame0[7][6] = 3'd0;
    frame0[7][7] = 3'd0;
    frame0[7][8] = 3'd0;
    frame0[7][9] = 3'd0;
    frame0[7][10] = 3'd0;
    frame0[7][11] = 3'd0;
    frame0[7][12] = 3'd1;
    frame0[7][13] = 3'd1;
    frame0[7][14] = 3'd3;
    frame0[7][15] = 3'd1;
    // frame0[7][16] = 3'd1;
    // frame0[7][17] = 3'd3;
    // frame0[7][18] = 3'd1;
    // frame0[7][19] = 3'd1;
    // frame0[7][20] = 3'd0;
    // frame0[7][21] = 3'd0;
    // frame0[7][22] = 3'd0;
    // frame0[7][23] = 3'd0;
    // frame0[7][24] = 3'd0;
    // frame0[7][25] = 3'd0;
    // frame0[7][26] = 3'd0;
    // frame0[7][27] = 3'd0;
    // frame0[7][28] = 3'd0;
    // frame0[7][29] = 3'd0;
    // frame0[7][30] = 3'd0;
    // frame0[7][31] = 3'd0;
    frame0[8][0] = 3'd0;
    frame0[8][1] = 3'd0;
    frame0[8][2] = 3'd0;
    frame0[8][3] = 3'd0;
    frame0[8][4] = 3'd0;
    frame0[8][5] = 3'd0;
    frame0[8][6] = 3'd0;
    frame0[8][7] = 3'd0;
    frame0[8][8] = 3'd0;
    frame0[8][9] = 3'd0;
    frame0[8][10] = 3'd0;
    frame0[8][11] = 3'd0;
    frame0[8][12] = 3'd0;
    frame0[8][13] = 3'd0;
    frame0[8][14] = 3'd1;
    frame0[8][15] = 3'd1;
    // frame0[8][16] = 3'd1;
    // frame0[8][17] = 3'd1;
    // frame0[8][18] = 3'd0;
    // frame0[8][19] = 3'd0;
    // frame0[8][20] = 3'd0;
    // frame0[8][21] = 3'd0;
    // frame0[8][22] = 3'd0;
    // frame0[8][23] = 3'd0;
    // frame0[8][24] = 3'd0;
    // frame0[8][25] = 3'd0;
    // frame0[8][26] = 3'd0;
    // frame0[8][27] = 3'd0;
    // frame0[8][28] = 3'd0;
    // frame0[8][29] = 3'd0;
    // frame0[8][30] = 3'd0;
    // frame0[8][31] = 3'd0;
    frame0[9][0] = 3'd0;
    frame0[9][1] = 3'd0;
    frame0[9][2] = 3'd0;
    frame0[9][3] = 3'd0;
    frame0[9][4] = 3'd0;
    frame0[9][5] = 3'd0;
    frame0[9][6] = 3'd0;
    frame0[9][7] = 3'd0;
    frame0[9][8] = 3'd0;
    frame0[9][9] = 3'd0;
    frame0[9][10] = 3'd0;
    frame0[9][11] = 3'd0;
    frame0[9][12] = 3'd0;
    frame0[9][13] = 3'd0;
    frame0[9][14] = 3'd1;
    frame0[9][15] = 3'd2;
    // frame0[9][16] = 3'd2;
    // frame0[9][17] = 3'd1;
    // frame0[9][18] = 3'd0;
    // frame0[9][19] = 3'd0;
    // frame0[9][20] = 3'd0;
    // frame0[9][21] = 3'd0;
    // frame0[9][22] = 3'd0;
    // frame0[9][23] = 3'd0;
    // frame0[9][24] = 3'd0;
    // frame0[9][25] = 3'd0;
    // frame0[9][26] = 3'd0;
    // frame0[9][27] = 3'd0;
    // frame0[9][28] = 3'd0;
    // frame0[9][29] = 3'd0;
    // frame0[9][30] = 3'd0;
    // frame0[9][31] = 3'd0;
    frame0[10][0] = 3'd0;
    frame0[10][1] = 3'd0;
    frame0[10][2] = 3'd0;
    frame0[10][3] = 3'd0;
    frame0[10][4] = 3'd0;
    frame0[10][5] = 3'd0;
    frame0[10][6] = 3'd0;
    frame0[10][7] = 3'd0;
    frame0[10][8] = 3'd0;
    frame0[10][9] = 3'd0;
    frame0[10][10] = 3'd0;
    frame0[10][11] = 3'd0;
    frame0[10][12] = 3'd0;
    frame0[10][13] = 3'd0;
    frame0[10][14] = 3'd1;
    frame0[10][15] = 3'd2;
    // frame0[10][16] = 3'd2;
    // frame0[10][17] = 3'd1;
    // frame0[10][18] = 3'd0;
    // frame0[10][19] = 3'd0;
    // frame0[10][20] = 3'd0;
    // frame0[10][21] = 3'd0;
    // frame0[10][22] = 3'd0;
    // frame0[10][23] = 3'd0;
    // frame0[10][24] = 3'd0;
    // frame0[10][25] = 3'd0;
    // frame0[10][26] = 3'd0;
    // frame0[10][27] = 3'd0;
    // frame0[10][28] = 3'd0;
    // frame0[10][29] = 3'd0;
    // frame0[10][30] = 3'd0;
    // frame0[10][31] = 3'd0;
    frame0[11][0] = 3'd0;
    frame0[11][1] = 3'd0;
    frame0[11][2] = 3'd0;
    frame0[11][3] = 3'd0;
    frame0[11][4] = 3'd0;
    frame0[11][5] = 3'd0;
    frame0[11][6] = 3'd0;
    frame0[11][7] = 3'd0;
    frame0[11][8] = 3'd0;
    frame0[11][9] = 3'd0;
    frame0[11][10] = 3'd0;
    frame0[11][11] = 3'd0;
    frame0[11][12] = 3'd0;
    frame0[11][13] = 3'd0;
    frame0[11][14] = 3'd1;
    frame0[11][15] = 3'd2;
    // frame0[11][16] = 3'd2;
    // frame0[11][17] = 3'd1;
    // frame0[11][18] = 3'd0;
    // frame0[11][19] = 3'd0;
    // frame0[11][20] = 3'd0;
    // frame0[11][21] = 3'd0;
    // frame0[11][22] = 3'd0;
    // frame0[11][23] = 3'd0;
    // frame0[11][24] = 3'd0;
    // frame0[11][25] = 3'd0;
    // frame0[11][26] = 3'd0;
    // frame0[11][27] = 3'd0;
    // frame0[11][28] = 3'd0;
    // frame0[11][29] = 3'd0;
    // frame0[11][30] = 3'd0;
    // frame0[11][31] = 3'd0;
    frame0[12][0] = 3'd0;
    frame0[12][1] = 3'd0;
    frame0[12][2] = 3'd0;
    frame0[12][3] = 3'd0;
    frame0[12][4] = 3'd0;
    frame0[12][5] = 3'd0;
    frame0[12][6] = 3'd0;
    frame0[12][7] = 3'd0;
    frame0[12][8] = 3'd0;
    frame0[12][9] = 3'd0;
    frame0[12][10] = 3'd0;
    frame0[12][11] = 3'd0;
    frame0[12][12] = 3'd0;
    frame0[12][13] = 3'd0;
    frame0[12][14] = 3'd1;
    frame0[12][15] = 3'd2;
    // frame0[12][16] = 3'd2;
    // frame0[12][17] = 3'd1;
    // frame0[12][18] = 3'd0;
    // frame0[12][19] = 3'd0;
    // frame0[12][20] = 3'd0;
    // frame0[12][21] = 3'd0;
    // frame0[12][22] = 3'd0;
    // frame0[12][23] = 3'd0;
    // frame0[12][24] = 3'd0;
    // frame0[12][25] = 3'd0;
    // frame0[12][26] = 3'd0;
    // frame0[12][27] = 3'd0;
    // frame0[12][28] = 3'd0;
    // frame0[12][29] = 3'd0;
    // frame0[12][30] = 3'd0;
    // frame0[12][31] = 3'd0;
    frame0[13][0] = 3'd0;
    frame0[13][1] = 3'd0;
    frame0[13][2] = 3'd0;
    frame0[13][3] = 3'd0;
    frame0[13][4] = 3'd0;
    frame0[13][5] = 3'd0;
    frame0[13][6] = 3'd0;
    frame0[13][7] = 3'd0;
    frame0[13][8] = 3'd0;
    frame0[13][9] = 3'd0;
    frame0[13][10] = 3'd0;
    frame0[13][11] = 3'd0;
    frame0[13][12] = 3'd0;
    frame0[13][13] = 3'd1;
    frame0[13][14] = 3'd1;
    frame0[13][15] = 3'd2;
    // frame0[13][16] = 3'd2;
    // frame0[13][17] = 3'd1;
    // frame0[13][18] = 3'd1;
    // frame0[13][19] = 3'd0;
    // frame0[13][20] = 3'd0;
    // frame0[13][21] = 3'd0;
    // frame0[13][22] = 3'd0;
    // frame0[13][23] = 3'd0;
    // frame0[13][24] = 3'd0;
    // frame0[13][25] = 3'd0;
    // frame0[13][26] = 3'd0;
    // frame0[13][27] = 3'd0;
    // frame0[13][28] = 3'd0;
    // frame0[13][29] = 3'd0;
    // frame0[13][30] = 3'd0;
    // frame0[13][31] = 3'd0;
    frame0[14][0] = 3'd0;
    frame0[14][1] = 3'd0;
    frame0[14][2] = 3'd0;
    frame0[14][3] = 3'd0;
    frame0[14][4] = 3'd0;
    frame0[14][5] = 3'd0;
    frame0[14][6] = 3'd0;
    frame0[14][7] = 3'd0;
    frame0[14][8] = 3'd0;
    frame0[14][9] = 3'd0;
    frame0[14][10] = 3'd0;
    frame0[14][11] = 3'd0;
    frame0[14][12] = 3'd1;
    frame0[14][13] = 3'd2;
    frame0[14][14] = 3'd4;
    frame0[14][15] = 3'd4;
    // frame0[14][16] = 3'd4;
    // frame0[14][17] = 3'd4;
    // frame0[14][18] = 3'd2;
    // frame0[14][19] = 3'd1;
    // frame0[14][20] = 3'd0;
    // frame0[14][21] = 3'd0;
    // frame0[14][22] = 3'd0;
    // frame0[14][23] = 3'd0;
    // frame0[14][24] = 3'd0;
    // frame0[14][25] = 3'd0;
    // frame0[14][26] = 3'd0;
    // frame0[14][27] = 3'd0;
    // frame0[14][28] = 3'd0;
    // frame0[14][29] = 3'd0;
    // frame0[14][30] = 3'd0;
    // frame0[14][31] = 3'd0;
    frame0[15][0] = 3'd0;
    frame0[15][1] = 3'd0;
    frame0[15][2] = 3'd0;
    frame0[15][3] = 3'd0;
    frame0[15][4] = 3'd0;
    frame0[15][5] = 3'd0;
    frame0[15][6] = 3'd0;
    frame0[15][7] = 3'd0;
    frame0[15][8] = 3'd0;
    frame0[15][9] = 3'd0;
    frame0[15][10] = 3'd0;
    frame0[15][11] = 3'd1;
    frame0[15][12] = 3'd2;
    frame0[15][13] = 3'd2;
    frame0[15][14] = 3'd4;
    frame0[15][15] = 3'd4;
    // frame0[15][16] = 3'd4;
    // frame0[15][17] = 3'd4;
    // frame0[15][18] = 3'd2;
    // frame0[15][19] = 3'd2;
    // frame0[15][20] = 3'd1;
    // frame0[15][21] = 3'd0;
    // frame0[15][22] = 3'd0;
    // frame0[15][23] = 3'd0;
    // frame0[15][24] = 3'd0;
    // frame0[15][25] = 3'd0;
    // frame0[15][26] = 3'd0;
    // frame0[15][27] = 3'd0;
    // frame0[15][28] = 3'd0;
    // frame0[15][29] = 3'd0;
    // frame0[15][30] = 3'd0;
    // frame0[15][31] = 3'd0;
    // frame0[16][0] = 3'd0;
    // frame0[16][1] = 3'd0;
    // frame0[16][2] = 3'd0;
    // frame0[16][3] = 3'd0;
    // frame0[16][4] = 3'd0;
    // frame0[16][5] = 3'd0;
    // frame0[16][6] = 3'd0;
    // frame0[16][7] = 3'd0;
    // frame0[16][8] = 3'd0;
    // frame0[16][9] = 3'd1;
    // frame0[16][10] = 3'd1;
    // frame0[16][11] = 3'd2;
    // frame0[16][12] = 3'd2;
    // frame0[16][13] = 3'd4;
    // frame0[16][14] = 3'd4;
    // frame0[16][15] = 3'd4;
    // frame0[16][16] = 3'd4;
    // frame0[16][17] = 3'd4;
    // frame0[16][18] = 3'd4;
    // frame0[16][19] = 3'd2;
    // frame0[16][20] = 3'd2;
    // frame0[16][21] = 3'd1;
    // frame0[16][22] = 3'd1;
    // frame0[16][23] = 3'd0;
    // frame0[16][24] = 3'd0;
    // frame0[16][25] = 3'd0;
    // frame0[16][26] = 3'd0;
    // frame0[16][27] = 3'd0;
    // frame0[16][28] = 3'd0;
    // frame0[16][29] = 3'd0;
    // frame0[16][30] = 3'd0;
    // frame0[16][31] = 3'd0;
    // frame0[17][0] = 3'd0;
    // frame0[17][1] = 3'd0;
    // frame0[17][2] = 3'd0;
    // frame0[17][3] = 3'd0;
    // frame0[17][4] = 3'd0;
    // frame0[17][5] = 3'd0;
    // frame0[17][6] = 3'd0;
    // frame0[17][7] = 3'd0;
    // frame0[17][8] = 3'd1;
    // frame0[17][9] = 3'd1;
    // frame0[17][10] = 3'd2;
    // frame0[17][11] = 3'd2;
    // frame0[17][12] = 3'd4;
    // frame0[17][13] = 3'd4;
    // frame0[17][14] = 3'd4;
    // frame0[17][15] = 3'd4;
    // frame0[17][16] = 3'd4;
    // frame0[17][17] = 3'd4;
    // frame0[17][18] = 3'd4;
    // frame0[17][19] = 3'd4;
    // frame0[17][20] = 3'd2;
    // frame0[17][21] = 3'd2;
    // frame0[17][22] = 3'd1;
    // frame0[17][23] = 3'd1;
    // frame0[17][24] = 3'd0;
    // frame0[17][25] = 3'd0;
    // frame0[17][26] = 3'd0;
    // frame0[17][27] = 3'd0;
    // frame0[17][28] = 3'd0;
    // frame0[17][29] = 3'd0;
    // frame0[17][30] = 3'd0;
    // frame0[17][31] = 3'd0;
    // frame0[18][0] = 3'd0;
    // frame0[18][1] = 3'd0;
    // frame0[18][2] = 3'd0;
    // frame0[18][3] = 3'd0;
    // frame0[18][4] = 3'd0;
    // frame0[18][5] = 3'd0;
    // frame0[18][6] = 3'd0;
    // frame0[18][7] = 3'd1;
    // frame0[18][8] = 3'd1;
    // frame0[18][9] = 3'd2;
    // frame0[18][10] = 3'd2;
    // frame0[18][11] = 3'd5;
    // frame0[18][12] = 3'd4;
    // frame0[18][13] = 3'd4;
    // frame0[18][14] = 3'd4;
    // frame0[18][15] = 3'd4;
    // frame0[18][16] = 3'd4;
    // frame0[18][17] = 3'd4;
    // frame0[18][18] = 3'd4;
    // frame0[18][19] = 3'd4;
    // frame0[18][20] = 3'd5;
    // frame0[18][21] = 3'd2;
    // frame0[18][22] = 3'd2;
    // frame0[18][23] = 3'd1;
    // frame0[18][24] = 3'd1;
    // frame0[18][25] = 3'd0;
    // frame0[18][26] = 3'd0;
    // frame0[18][27] = 3'd0;
    // frame0[18][28] = 3'd0;
    // frame0[18][29] = 3'd0;
    // frame0[18][30] = 3'd0;
    // frame0[18][31] = 3'd0;
    // frame0[19][0] = 3'd0;
    // frame0[19][1] = 3'd0;
    // frame0[19][2] = 3'd0;
    // frame0[19][3] = 3'd0;
    // frame0[19][4] = 3'd0;
    // frame0[19][5] = 3'd0;
    // frame0[19][6] = 3'd0;
    // frame0[19][7] = 3'd1;
    // frame0[19][8] = 3'd2;
    // frame0[19][9] = 3'd2;
    // frame0[19][10] = 3'd2;
    // frame0[19][11] = 3'd5;
    // frame0[19][12] = 3'd4;
    // frame0[19][13] = 3'd4;
    // frame0[19][14] = 3'd4;
    // frame0[19][15] = 3'd4;
    // frame0[19][16] = 3'd4;
    // frame0[19][17] = 3'd4;
    // frame0[19][18] = 3'd4;
    // frame0[19][19] = 3'd4;
    // frame0[19][20] = 3'd5;
    // frame0[19][21] = 3'd2;
    // frame0[19][22] = 3'd2;
    // frame0[19][23] = 3'd2;
    // frame0[19][24] = 3'd1;
    // frame0[19][25] = 3'd0;
    // frame0[19][26] = 3'd0;
    // frame0[19][27] = 3'd0;
    // frame0[19][28] = 3'd0;
    // frame0[19][29] = 3'd0;
    // frame0[19][30] = 3'd0;
    // frame0[19][31] = 3'd0;
    // frame0[20][0] = 3'd0;
    // frame0[20][1] = 3'd0;
    // frame0[20][2] = 3'd0;
    // frame0[20][3] = 3'd0;
    // frame0[20][4] = 3'd0;
    // frame0[20][5] = 3'd0;
    // frame0[20][6] = 3'd0;
    // frame0[20][7] = 3'd1;
    // frame0[20][8] = 3'd2;
    // frame0[20][9] = 3'd2;
    // frame0[20][10] = 3'd1;
    // frame0[20][11] = 3'd5;
    // frame0[20][12] = 3'd4;
    // frame0[20][13] = 3'd4;
    // frame0[20][14] = 3'd4;
    // frame0[20][15] = 3'd4;
    // frame0[20][16] = 3'd4;
    // frame0[20][17] = 3'd4;
    // frame0[20][18] = 3'd4;
    // frame0[20][19] = 3'd4;
    // frame0[20][20] = 3'd5;
    // frame0[20][21] = 3'd1;
    // frame0[20][22] = 3'd2;
    // frame0[20][23] = 3'd2;
    // frame0[20][24] = 3'd1;
    // frame0[20][25] = 3'd0;
    // frame0[20][26] = 3'd0;
    // frame0[20][27] = 3'd0;
    // frame0[20][28] = 3'd0;
    // frame0[20][29] = 3'd0;
    // frame0[20][30] = 3'd0;
    // frame0[20][31] = 3'd0;
    // frame0[21][0] = 3'd0;
    // frame0[21][1] = 3'd0;
    // frame0[21][2] = 3'd0;
    // frame0[21][3] = 3'd0;
    // frame0[21][4] = 3'd0;
    // frame0[21][5] = 3'd0;
    // frame0[21][6] = 3'd0;
    // frame0[21][7] = 3'd1;
    // frame0[21][8] = 3'd1;
    // frame0[21][9] = 3'd2;
    // frame0[21][10] = 3'd1;
    // frame0[21][11] = 3'd2;
    // frame0[21][12] = 3'd5;
    // frame0[21][13] = 3'd4;
    // frame0[21][14] = 3'd4;
    // frame0[21][15] = 3'd4;
    // frame0[21][16] = 3'd4;
    // frame0[21][17] = 3'd4;
    // frame0[21][18] = 3'd4;
    // frame0[21][19] = 3'd5;
    // frame0[21][20] = 3'd2;
    // frame0[21][21] = 3'd1;
    // frame0[21][22] = 3'd2;
    // frame0[21][23] = 3'd1;
    // frame0[21][24] = 3'd1;
    // frame0[21][25] = 3'd0;
    // frame0[21][26] = 3'd0;
    // frame0[21][27] = 3'd0;
    // frame0[21][28] = 3'd0;
    // frame0[21][29] = 3'd0;
    // frame0[21][30] = 3'd0;
    // frame0[21][31] = 3'd0;
    // frame0[22][0] = 3'd0;
    // frame0[22][1] = 3'd0;
    // frame0[22][2] = 3'd0;
    // frame0[22][3] = 3'd0;
    // frame0[22][4] = 3'd0;
    // frame0[22][5] = 3'd0;
    // frame0[22][6] = 3'd0;
    // frame0[22][7] = 3'd0;
    // frame0[22][8] = 3'd1;
    // frame0[22][9] = 3'd1;
    // frame0[22][10] = 3'd1;
    // frame0[22][11] = 3'd2;
    // frame0[22][12] = 3'd2;
    // frame0[22][13] = 3'd5;
    // frame0[22][14] = 3'd4;
    // frame0[22][15] = 3'd4;
    // frame0[22][16] = 3'd4;
    // frame0[22][17] = 3'd4;
    // frame0[22][18] = 3'd5;
    // frame0[22][19] = 3'd2;
    // frame0[22][20] = 3'd2;
    // frame0[22][21] = 3'd1;
    // frame0[22][22] = 3'd1;
    // frame0[22][23] = 3'd1;
    // frame0[22][24] = 3'd0;
    // frame0[22][25] = 3'd0;
    // frame0[22][26] = 3'd0;
    // frame0[22][27] = 3'd0;
    // frame0[22][28] = 3'd0;
    // frame0[22][29] = 3'd0;
    // frame0[22][30] = 3'd0;
    // frame0[22][31] = 3'd0;
    // frame0[23][0] = 3'd0;
    // frame0[23][1] = 3'd0;
    // frame0[23][2] = 3'd0;
    // frame0[23][3] = 3'd0;
    // frame0[23][4] = 3'd0;
    // frame0[23][5] = 3'd0;
    // frame0[23][6] = 3'd0;
    // frame0[23][7] = 3'd0;
    // frame0[23][8] = 3'd0;
    // frame0[23][9] = 3'd1;
    // frame0[23][10] = 3'd1;
    // frame0[23][11] = 3'd1;
    // frame0[23][12] = 3'd2;
    // frame0[23][13] = 3'd2;
    // frame0[23][14] = 3'd5;
    // frame0[23][15] = 3'd5;
    // frame0[23][16] = 3'd5;
    // frame0[23][17] = 3'd5;
    // frame0[23][18] = 3'd2;
    // frame0[23][19] = 3'd2;
    // frame0[23][20] = 3'd1;
    // frame0[23][21] = 3'd1;
    // frame0[23][22] = 3'd1;
    // frame0[23][23] = 3'd0;
    // frame0[23][24] = 3'd0;
    // frame0[23][25] = 3'd0;
    // frame0[23][26] = 3'd0;
    // frame0[23][27] = 3'd0;
    // frame0[23][28] = 3'd0;
    // frame0[23][29] = 3'd0;
    // frame0[23][30] = 3'd0;
    // frame0[23][31] = 3'd0;
    // frame0[24][0] = 3'd0;
    // frame0[24][1] = 3'd0;
    // frame0[24][2] = 3'd0;
    // frame0[24][3] = 3'd0;
    // frame0[24][4] = 3'd0;
    // frame0[24][5] = 3'd0;
    // frame0[24][6] = 3'd0;
    // frame0[24][7] = 3'd0;
    // frame0[24][8] = 3'd0;
    // frame0[24][9] = 3'd0;
    // frame0[24][10] = 3'd0;
    // frame0[24][11] = 3'd1;
    // frame0[24][12] = 3'd1;
    // frame0[24][13] = 3'd2;
    // frame0[24][14] = 3'd2;
    // frame0[24][15] = 3'd5;
    // frame0[24][16] = 3'd5;
    // frame0[24][17] = 3'd2;
    // frame0[24][18] = 3'd2;
    // frame0[24][19] = 3'd1;
    // frame0[24][20] = 3'd1;
    // frame0[24][21] = 3'd0;
    // frame0[24][22] = 3'd0;
    // frame0[24][23] = 3'd0;
    // frame0[24][24] = 3'd0;
    // frame0[24][25] = 3'd0;
    // frame0[24][26] = 3'd0;
    // frame0[24][27] = 3'd0;
    // frame0[24][28] = 3'd0;
    // frame0[24][29] = 3'd0;
    // frame0[24][30] = 3'd0;
    // frame0[24][31] = 3'd0;
    // frame0[25][0] = 3'd0;
    // frame0[25][1] = 3'd0;
    // frame0[25][2] = 3'd0;
    // frame0[25][3] = 3'd0;
    // frame0[25][4] = 3'd0;
    // frame0[25][5] = 3'd0;
    // frame0[25][6] = 3'd0;
    // frame0[25][7] = 3'd0;
    // frame0[25][8] = 3'd0;
    // frame0[25][9] = 3'd0;
    // frame0[25][10] = 3'd0;
    // frame0[25][11] = 3'd0;
    // frame0[25][12] = 3'd1;
    // frame0[25][13] = 3'd1;
    // frame0[25][14] = 3'd2;
    // frame0[25][15] = 3'd2;
    // frame0[25][16] = 3'd2;
    // frame0[25][17] = 3'd2;
    // frame0[25][18] = 3'd1;
    // frame0[25][19] = 3'd1;
    // frame0[25][20] = 3'd0;
    // frame0[25][21] = 3'd0;
    // frame0[25][22] = 3'd0;
    // frame0[25][23] = 3'd0;
    // frame0[25][24] = 3'd0;
    // frame0[25][25] = 3'd0;
    // frame0[25][26] = 3'd0;
    // frame0[25][27] = 3'd0;
    // frame0[25][28] = 3'd0;
    // frame0[25][29] = 3'd0;
    // frame0[25][30] = 3'd0;
    // frame0[25][31] = 3'd0;
    // frame0[26][0] = 3'd0;
    // frame0[26][1] = 3'd0;
    // frame0[26][2] = 3'd0;
    // frame0[26][3] = 3'd0;
    // frame0[26][4] = 3'd0;
    // frame0[26][5] = 3'd0;
    // frame0[26][6] = 3'd0;
    // frame0[26][7] = 3'd0;
    // frame0[26][8] = 3'd0;
    // frame0[26][9] = 3'd0;
    // frame0[26][10] = 3'd0;
    // frame0[26][11] = 3'd0;
    // frame0[26][12] = 3'd1;
    // frame0[26][13] = 3'd0;
    // frame0[26][14] = 3'd1;
    // frame0[26][15] = 3'd2;
    // frame0[26][16] = 3'd2;
    // frame0[26][17] = 3'd1;
    // frame0[26][18] = 3'd0;
    // frame0[26][19] = 3'd1;
    // frame0[26][20] = 3'd0;
    // frame0[26][21] = 3'd0;
    // frame0[26][22] = 3'd0;
    // frame0[26][23] = 3'd0;
    // frame0[26][24] = 3'd0;
    // frame0[26][25] = 3'd0;
    // frame0[26][26] = 3'd0;
    // frame0[26][27] = 3'd0;
    // frame0[26][28] = 3'd0;
    // frame0[26][29] = 3'd0;
    // frame0[26][30] = 3'd0;
    // frame0[26][31] = 3'd0;
    // frame0[27][0] = 3'd0;
    // frame0[27][1] = 3'd0;
    // frame0[27][2] = 3'd0;
    // frame0[27][3] = 3'd0;
    // frame0[27][4] = 3'd0;
    // frame0[27][5] = 3'd0;
    // frame0[27][6] = 3'd0;
    // frame0[27][7] = 3'd0;
    // frame0[27][8] = 3'd0;
    // frame0[27][9] = 3'd0;
    // frame0[27][10] = 3'd0;
    // frame0[27][11] = 3'd0;
    // frame0[27][12] = 3'd1;
    // frame0[27][13] = 3'd0;
    // frame0[27][14] = 3'd0;
    // frame0[27][15] = 3'd1;
    // frame0[27][16] = 3'd1;
    // frame0[27][17] = 3'd0;
    // frame0[27][18] = 3'd0;
    // frame0[27][19] = 3'd1;
    // frame0[27][20] = 3'd0;
    // frame0[27][21] = 3'd0;
    // frame0[27][22] = 3'd0;
    // frame0[27][23] = 3'd0;
    // frame0[27][24] = 3'd0;
    // frame0[27][25] = 3'd0;
    // frame0[27][26] = 3'd0;
    // frame0[27][27] = 3'd0;
    // frame0[27][28] = 3'd0;
    // frame0[27][29] = 3'd0;
    // frame0[27][30] = 3'd0;
    // frame0[27][31] = 3'd0;
    // frame0[28][0] = 3'd0;
    // frame0[28][1] = 3'd0;
    // frame0[28][2] = 3'd0;
    // frame0[28][3] = 3'd0;
    // frame0[28][4] = 3'd0;
    // frame0[28][5] = 3'd0;
    // frame0[28][6] = 3'd0;
    // frame0[28][7] = 3'd0;
    // frame0[28][8] = 3'd0;
    // frame0[28][9] = 3'd0;
    // frame0[28][10] = 3'd0;
    // frame0[28][11] = 3'd0;
    // frame0[28][12] = 3'd1;
    // frame0[28][13] = 3'd0;
    // frame0[28][14] = 3'd0;
    // frame0[28][15] = 3'd0;
    // frame0[28][16] = 3'd0;
    // frame0[28][17] = 3'd0;
    // frame0[28][18] = 3'd0;
    // frame0[28][19] = 3'd1;
    // frame0[28][20] = 3'd0;
    // frame0[28][21] = 3'd0;
    // frame0[28][22] = 3'd0;
    // frame0[28][23] = 3'd0;
    // frame0[28][24] = 3'd0;
    // frame0[28][25] = 3'd0;
    // frame0[28][26] = 3'd0;
    // frame0[28][27] = 3'd0;
    // frame0[28][28] = 3'd0;
    // frame0[28][29] = 3'd0;
    // frame0[28][30] = 3'd0;
    // frame0[28][31] = 3'd0;
    // frame0[29][0] = 3'd0;
    // frame0[29][1] = 3'd0;
    // frame0[29][2] = 3'd0;
    // frame0[29][3] = 3'd0;
    // frame0[29][4] = 3'd0;
    // frame0[29][5] = 3'd0;
    // frame0[29][6] = 3'd0;
    // frame0[29][7] = 3'd0;
    // frame0[29][8] = 3'd0;
    // frame0[29][9] = 3'd0;
    // frame0[29][10] = 3'd0;
    // frame0[29][11] = 3'd0;
    // frame0[29][12] = 3'd1;
    // frame0[29][13] = 3'd0;
    // frame0[29][14] = 3'd0;
    // frame0[29][15] = 3'd0;
    // frame0[29][16] = 3'd0;
    // frame0[29][17] = 3'd0;
    // frame0[29][18] = 3'd0;
    // frame0[29][19] = 3'd1;
    // frame0[29][20] = 3'd0;
    // frame0[29][21] = 3'd0;
    // frame0[29][22] = 3'd0;
    // frame0[29][23] = 3'd0;
    // frame0[29][24] = 3'd0;
    // frame0[29][25] = 3'd0;
    // frame0[29][26] = 3'd0;
    // frame0[29][27] = 3'd0;
    // frame0[29][28] = 3'd0;
    // frame0[29][29] = 3'd0;
    // frame0[29][30] = 3'd0;
    // frame0[29][31] = 3'd0;
    // frame0[30][0] = 3'd0;
    // frame0[30][1] = 3'd0;
    // frame0[30][2] = 3'd0;
    // frame0[30][3] = 3'd0;
    // frame0[30][4] = 3'd0;
    // frame0[30][5] = 3'd0;
    // frame0[30][6] = 3'd0;
    // frame0[30][7] = 3'd0;
    // frame0[30][8] = 3'd0;
    // frame0[30][9] = 3'd0;
    // frame0[30][10] = 3'd0;
    // frame0[30][11] = 3'd1;
    // frame0[30][12] = 3'd1;
    // frame0[30][13] = 3'd1;
    // frame0[30][14] = 3'd0;
    // frame0[30][15] = 3'd0;
    // frame0[30][16] = 3'd0;
    // frame0[30][17] = 3'd0;
    // frame0[30][18] = 3'd1;
    // frame0[30][19] = 3'd1;
    // frame0[30][20] = 3'd1;
    // frame0[30][21] = 3'd0;
    // frame0[30][22] = 3'd0;
    // frame0[30][23] = 3'd0;
    // frame0[30][24] = 3'd0;
    // frame0[30][25] = 3'd0;
    // frame0[30][26] = 3'd0;
    // frame0[30][27] = 3'd0;
    // frame0[30][28] = 3'd0;
    // frame0[30][29] = 3'd0;
    // frame0[30][30] = 3'd0;
    // frame0[30][31] = 3'd0;
    // frame0[31][0] = 3'd0;
    // frame0[31][1] = 3'd0;
    // frame0[31][2] = 3'd0;
    // frame0[31][3] = 3'd0;
    // frame0[31][4] = 3'd0;
    // frame0[31][5] = 3'd0;
    // frame0[31][6] = 3'd0;
    // frame0[31][7] = 3'd0;
    // frame0[31][8] = 3'd0;
    // frame0[31][9] = 3'd0;
    // frame0[31][10] = 3'd1;
    // frame0[31][11] = 3'd0;
    // frame0[31][12] = 3'd1;
    // frame0[31][13] = 3'd0;
    // frame0[31][14] = 3'd1;
    // frame0[31][15] = 3'd0;
    // frame0[31][16] = 3'd0;
    // frame0[31][17] = 3'd1;
    // frame0[31][18] = 3'd0;
    // frame0[31][19] = 3'd1;
    // frame0[31][20] = 3'd0;
    // frame0[31][21] = 3'd1;
    // frame0[31][22] = 3'd0;
    // frame0[31][23] = 3'd0;
    // frame0[31][24] = 3'd0;
    // frame0[31][25] = 3'd0;
    // frame0[31][26] = 3'd0;
    // frame0[31][27] = 3'd0;
    // frame0[31][28] = 3'd0;
    // frame0[31][29] = 3'd0;
    // frame0[31][30] = 3'd0;
    // frame0[31][31] = 3'd0;
end